VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Burrows_Katie
  CLASS BLOCK ;
  FOREIGN tt_um_Burrows_Katie ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 57.065 54.275 57.075 54.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 210.765 42.820 212.650 45.305 ;
    END
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END VPWR
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 17.639999 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.410000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.410000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.095000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER pwell ;
        RECT 52.645 212.180 53.315 212.260 ;
        RECT 52.645 209.390 58.585 212.180 ;
      LAYER nwell ;
        RECT 98.120 210.370 104.540 215.650 ;
        RECT 106.200 210.370 112.620 215.650 ;
      LAYER pwell ;
        RECT 52.645 209.310 53.315 209.390 ;
        RECT 52.645 207.480 53.315 207.560 ;
        RECT 52.645 204.690 58.585 207.480 ;
      LAYER nwell ;
        RECT 63.305 206.300 65.725 209.580 ;
        RECT 92.285 206.335 94.705 209.615 ;
      LAYER pwell ;
        RECT 52.645 204.610 53.315 204.690 ;
      LAYER nwell ;
        RECT 98.120 203.380 104.540 208.660 ;
        RECT 106.200 203.380 112.620 208.660 ;
      LAYER pwell ;
        RECT 52.645 200.945 53.315 201.025 ;
        RECT 52.645 198.155 58.585 200.945 ;
        RECT 52.645 198.075 53.315 198.155 ;
      LAYER nwell ;
        RECT 76.830 196.990 83.250 202.270 ;
        RECT 98.120 196.390 104.540 201.670 ;
        RECT 106.200 196.390 112.620 201.670 ;
      LAYER pwell ;
        RECT 52.645 196.135 53.315 196.215 ;
        RECT 52.645 193.345 58.585 196.135 ;
        RECT 52.645 193.265 53.315 193.345 ;
      LAYER nwell ;
        RECT 76.830 190.075 83.250 195.355 ;
        RECT 98.120 189.365 104.540 194.645 ;
        RECT 106.200 189.365 112.620 194.645 ;
      LAYER pwell ;
        RECT 45.550 187.740 46.220 187.820 ;
        RECT 45.550 184.950 53.490 187.740 ;
        RECT 45.550 184.870 46.220 184.950 ;
        RECT 45.550 183.265 46.220 183.345 ;
        RECT 45.550 180.475 53.490 183.265 ;
        RECT 45.550 180.395 46.220 180.475 ;
        RECT 45.550 178.650 46.220 178.730 ;
        RECT 45.550 175.860 53.490 178.650 ;
        RECT 45.550 175.780 46.220 175.860 ;
        RECT 45.530 173.075 46.200 173.155 ;
        RECT 45.530 170.285 53.470 173.075 ;
      LAYER nwell ;
        RECT 88.680 172.365 91.100 175.645 ;
        RECT 106.425 170.750 112.845 176.030 ;
      LAYER pwell ;
        RECT 45.530 170.205 46.200 170.285 ;
        RECT 45.530 168.560 46.200 168.640 ;
        RECT 45.530 165.770 53.470 168.560 ;
        RECT 45.530 165.690 46.200 165.770 ;
        RECT 45.530 163.970 46.200 164.050 ;
        RECT 45.530 161.180 53.470 163.970 ;
      LAYER nwell ;
        RECT 88.675 162.365 91.095 165.645 ;
        RECT 106.425 163.640 112.845 168.920 ;
      LAYER pwell ;
        RECT 45.530 161.100 46.200 161.180 ;
        RECT 43.430 107.225 44.100 107.305 ;
        RECT 43.430 102.435 49.370 107.225 ;
        RECT 43.430 102.355 44.100 102.435 ;
      LAYER nwell ;
        RECT 52.695 102.245 59.115 107.525 ;
        RECT 62.845 102.245 69.265 107.525 ;
        RECT 72.125 102.200 78.545 107.480 ;
      LAYER pwell ;
        RECT 43.430 97.410 44.100 97.490 ;
        RECT 43.430 92.620 49.370 97.410 ;
        RECT 43.430 92.540 44.100 92.620 ;
      LAYER nwell ;
        RECT 52.695 92.350 59.115 97.630 ;
        RECT 62.845 92.370 69.265 97.650 ;
        RECT 72.125 92.310 78.545 97.590 ;
      LAYER pwell ;
        RECT 43.430 87.250 44.100 87.330 ;
        RECT 43.430 82.460 49.370 87.250 ;
        RECT 43.430 82.380 44.100 82.460 ;
      LAYER nwell ;
        RECT 52.695 82.305 59.115 87.585 ;
        RECT 62.845 82.430 69.265 87.710 ;
        RECT 72.080 82.475 78.500 87.755 ;
        RECT 95.525 81.215 101.945 94.185 ;
        RECT 113.870 81.215 120.290 94.185 ;
      LAYER pwell ;
        RECT 43.430 78.185 44.100 78.265 ;
        RECT 43.430 73.395 49.370 78.185 ;
        RECT 43.430 73.315 44.100 73.395 ;
      LAYER nwell ;
        RECT 52.695 73.105 59.115 78.385 ;
        RECT 62.845 73.010 69.265 78.290 ;
        RECT 72.125 72.915 78.545 78.195 ;
      LAYER pwell ;
        RECT 49.115 69.970 49.785 70.050 ;
        RECT 49.115 66.180 56.055 69.970 ;
        RECT 49.115 66.100 49.785 66.180 ;
        RECT 49.115 63.280 49.785 63.360 ;
        RECT 49.115 59.490 56.055 63.280 ;
        RECT 49.115 59.410 49.785 59.490 ;
        RECT 49.115 56.590 49.785 56.670 ;
        RECT 49.115 52.800 56.055 56.590 ;
      LAYER nwell ;
        RECT 62.040 54.450 70.460 68.190 ;
        RECT 74.395 54.870 82.815 68.670 ;
        RECT 95.220 62.925 101.640 75.895 ;
        RECT 113.875 62.680 120.295 75.650 ;
      LAYER pwell ;
        RECT 49.115 52.720 49.785 52.800 ;
        RECT 49.115 49.950 49.785 50.030 ;
        RECT 49.115 46.160 56.055 49.950 ;
        RECT 49.115 46.080 49.785 46.160 ;
        RECT 35.645 43.750 36.315 43.830 ;
        RECT 45.770 43.750 46.440 43.830 ;
        RECT 35.645 39.960 42.685 43.750 ;
        RECT 45.770 39.960 52.810 43.750 ;
        RECT 35.645 39.880 36.315 39.960 ;
        RECT 45.770 39.880 46.440 39.960 ;
      LAYER nwell ;
        RECT 62.295 37.745 70.715 51.485 ;
        RECT 74.415 37.225 82.835 51.025 ;
        RECT 111.060 43.650 119.480 55.990 ;
      LAYER pwell ;
        RECT 35.645 37.055 36.315 37.135 ;
        RECT 45.770 37.055 46.440 37.135 ;
        RECT 35.645 33.265 42.685 37.055 ;
        RECT 45.770 33.265 52.810 37.055 ;
        RECT 70.125 34.295 70.795 34.375 ;
        RECT 56.675 34.120 57.345 34.200 ;
        RECT 35.645 33.185 36.315 33.265 ;
        RECT 45.770 33.185 46.440 33.265 ;
        RECT 56.675 32.700 64.615 34.120 ;
        RECT 70.125 32.875 78.065 34.295 ;
        RECT 70.125 32.795 70.795 32.875 ;
        RECT 56.675 32.620 57.345 32.700 ;
        RECT 35.645 30.940 36.315 31.020 ;
        RECT 45.770 30.940 46.440 31.020 ;
        RECT 35.645 27.150 42.685 30.940 ;
        RECT 45.770 27.150 52.810 30.940 ;
        RECT 35.645 27.070 36.315 27.150 ;
        RECT 45.770 27.070 46.440 27.150 ;
        RECT 35.645 24.535 36.315 24.615 ;
        RECT 45.770 24.535 46.440 24.615 ;
        RECT 35.645 20.745 42.685 24.535 ;
        RECT 45.770 20.745 52.810 24.535 ;
        RECT 35.645 20.665 36.315 20.745 ;
        RECT 45.770 20.665 46.440 20.745 ;
      LAYER li1 ;
        RECT 98.995 215.630 99.525 216.160 ;
        RECT 107.275 215.630 107.805 216.160 ;
        RECT 99.110 215.235 99.410 215.630 ;
        RECT 98.805 215.065 103.555 215.235 ;
        RECT 103.990 214.570 104.320 215.315 ;
        RECT 107.390 215.235 107.690 215.630 ;
        RECT 106.885 215.065 111.635 215.235 ;
        RECT 104.605 214.570 105.135 214.705 ;
        RECT 103.990 214.240 105.135 214.570 ;
        RECT 52.815 211.265 53.145 212.090 ;
        RECT 53.850 212.010 54.550 213.200 ;
        RECT 97.600 212.970 98.200 213.570 ;
        RECT 53.580 211.840 58.330 212.010 ;
        RECT 51.905 210.565 53.145 211.265 ;
        RECT 52.815 209.480 53.145 210.565 ;
        RECT 59.010 210.420 59.540 210.950 ;
        RECT 98.805 210.785 103.555 210.955 ;
        RECT 103.240 210.370 103.410 210.785 ;
        RECT 103.990 210.705 104.320 214.240 ;
        RECT 104.605 214.175 105.135 214.240 ;
        RECT 112.070 214.415 112.400 215.315 ;
        RECT 112.705 214.415 113.235 214.555 ;
        RECT 112.070 214.085 113.235 214.415 ;
        RECT 105.795 213.110 106.395 213.710 ;
        RECT 106.885 210.785 111.635 210.955 ;
        RECT 107.090 210.640 107.395 210.785 ;
        RECT 112.070 210.705 112.400 214.085 ;
        RECT 112.705 214.025 113.235 214.085 ;
        RECT 107.095 210.370 107.395 210.640 ;
        RECT 53.580 209.560 58.330 209.730 ;
        RECT 64.110 209.630 64.640 210.160 ;
        RECT 93.195 209.630 93.725 210.160 ;
        RECT 103.060 209.840 103.590 210.370 ;
        RECT 106.980 209.840 107.510 210.370 ;
        RECT 53.650 209.230 53.950 209.560 ;
        RECT 53.535 208.700 54.065 209.230 ;
        RECT 64.225 209.165 64.395 209.630 ;
        RECT 65.195 209.245 65.525 209.265 ;
        RECT 64.030 208.995 64.700 209.165 ;
        RECT 52.815 206.365 53.145 207.390 ;
        RECT 53.840 207.310 54.540 208.135 ;
        RECT 62.570 207.920 63.460 208.810 ;
        RECT 53.580 207.140 58.330 207.310 ;
        RECT 64.030 206.820 64.700 206.885 ;
        RECT 51.905 205.665 53.145 206.365 ;
        RECT 64.015 206.715 64.700 206.820 ;
        RECT 64.015 206.355 64.415 206.715 ;
        RECT 65.175 206.635 65.525 209.245 ;
        RECT 93.320 209.200 93.620 209.630 ;
        RECT 93.010 209.030 93.680 209.200 ;
        RECT 93.320 208.995 93.620 209.030 ;
        RECT 91.480 207.920 92.370 208.810 ;
        RECT 93.010 206.750 93.680 206.920 ;
        RECT 94.155 206.810 94.485 209.280 ;
        RECT 98.995 208.435 99.525 208.965 ;
        RECT 107.275 208.435 107.805 208.965 ;
        RECT 99.110 208.245 99.410 208.435 ;
        RECT 98.805 208.075 103.555 208.245 ;
        RECT 59.010 205.765 59.540 206.295 ;
        RECT 63.930 205.825 64.460 206.355 ;
        RECT 52.815 204.780 53.145 205.665 ;
        RECT 65.195 205.280 65.525 206.635 ;
        RECT 93.320 206.375 93.620 206.750 ;
        RECT 94.130 206.670 94.485 206.810 ;
        RECT 103.990 207.650 104.320 208.325 ;
        RECT 107.390 208.245 107.690 208.435 ;
        RECT 106.885 208.075 111.635 208.245 ;
        RECT 104.625 207.650 105.155 207.790 ;
        RECT 103.990 207.320 105.155 207.650 ;
        RECT 93.195 205.845 93.725 206.375 ;
        RECT 94.130 205.375 94.460 206.670 ;
        RECT 97.600 205.795 98.200 206.395 ;
        RECT 53.580 204.860 58.330 205.030 ;
        RECT 53.610 204.420 53.910 204.860 ;
        RECT 65.195 204.850 65.735 205.280 ;
        RECT 65.205 204.750 65.735 204.850 ;
        RECT 94.005 204.845 94.535 205.375 ;
        RECT 53.495 203.890 54.025 204.420 ;
        RECT 98.805 203.795 103.555 203.965 ;
        RECT 103.325 203.305 103.495 203.795 ;
        RECT 103.990 203.715 104.320 207.320 ;
        RECT 104.625 207.260 105.155 207.320 ;
        RECT 112.070 207.650 112.400 208.325 ;
        RECT 112.705 207.650 113.235 207.790 ;
        RECT 112.070 207.320 113.235 207.650 ;
        RECT 105.795 206.030 106.395 206.630 ;
        RECT 106.885 203.795 111.635 203.965 ;
        RECT 107.180 203.305 107.480 203.795 ;
        RECT 112.070 203.715 112.400 207.320 ;
        RECT 112.705 207.260 113.235 207.320 ;
        RECT 81.475 201.855 82.175 203.075 ;
        RECT 103.145 202.775 103.675 203.305 ;
        RECT 107.065 202.775 107.595 203.305 ;
        RECT 52.815 199.830 53.145 200.855 ;
        RECT 53.765 200.775 54.465 201.705 ;
        RECT 77.515 201.685 82.265 201.855 ;
        RECT 82.700 201.815 83.030 201.935 ;
        RECT 82.700 201.115 84.000 201.815 ;
        RECT 98.995 201.460 99.525 201.990 ;
        RECT 107.275 201.530 107.805 202.060 ;
        RECT 99.110 201.255 99.410 201.460 ;
        RECT 53.580 200.605 58.330 200.775 ;
        RECT 51.905 199.130 53.145 199.830 ;
        RECT 59.010 199.370 59.540 199.900 ;
        RECT 76.275 199.385 76.805 199.915 ;
        RECT 52.815 198.245 53.145 199.130 ;
        RECT 53.580 198.325 58.330 198.495 ;
        RECT 53.665 198.000 53.965 198.325 ;
        RECT 53.550 197.470 54.080 198.000 ;
        RECT 77.515 197.405 82.265 197.575 ;
        RECT 77.835 197.020 78.135 197.405 ;
        RECT 82.700 197.325 83.030 201.115 ;
        RECT 98.805 201.085 103.555 201.255 ;
        RECT 103.990 200.475 104.320 201.335 ;
        RECT 107.390 201.255 107.690 201.530 ;
        RECT 106.885 201.085 111.635 201.255 ;
        RECT 104.625 200.475 105.155 200.680 ;
        RECT 103.990 200.150 105.155 200.475 ;
        RECT 112.070 200.475 112.400 201.335 ;
        RECT 112.705 200.475 113.235 200.680 ;
        RECT 112.070 200.150 113.235 200.475 ;
        RECT 103.990 200.145 105.055 200.150 ;
        RECT 112.070 200.145 113.135 200.150 ;
        RECT 97.600 198.845 98.200 199.445 ;
        RECT 52.815 195.140 53.145 196.045 ;
        RECT 53.820 195.965 54.520 196.780 ;
        RECT 77.720 196.490 78.250 197.020 ;
        RECT 98.805 196.805 103.555 196.975 ;
        RECT 103.325 196.425 103.495 196.805 ;
        RECT 103.990 196.725 104.320 200.145 ;
        RECT 105.795 199.160 106.395 199.760 ;
        RECT 106.885 196.805 111.635 196.975 ;
        RECT 107.180 196.425 107.480 196.805 ;
        RECT 112.070 196.725 112.400 200.145 ;
        RECT 53.580 195.795 58.330 195.965 ;
        RECT 51.905 194.440 53.145 195.140 ;
        RECT 81.475 194.940 82.175 195.970 ;
        RECT 103.145 195.895 103.675 196.425 ;
        RECT 107.065 195.895 107.595 196.425 ;
        RECT 52.815 193.435 53.145 194.440 ;
        RECT 59.010 194.325 59.540 194.855 ;
        RECT 77.515 194.770 82.265 194.940 ;
        RECT 82.700 194.920 83.030 195.020 ;
        RECT 82.700 194.220 84.000 194.920 ;
        RECT 98.995 194.485 99.525 195.015 ;
        RECT 107.275 194.550 107.805 195.080 ;
        RECT 99.175 194.230 99.345 194.485 ;
        RECT 53.580 193.515 58.330 193.685 ;
        RECT 53.630 193.180 53.930 193.515 ;
        RECT 53.550 192.650 54.080 193.180 ;
        RECT 76.255 192.110 76.785 192.640 ;
        RECT 77.515 190.490 82.265 190.660 ;
        RECT 77.835 190.155 78.135 190.490 ;
        RECT 82.700 190.410 83.030 194.220 ;
        RECT 98.805 194.060 103.555 194.230 ;
        RECT 103.990 193.375 104.320 194.310 ;
        RECT 107.390 194.230 107.690 194.550 ;
        RECT 106.885 194.060 111.635 194.230 ;
        RECT 104.625 193.375 105.155 193.615 ;
        RECT 103.990 193.085 105.155 193.375 ;
        RECT 103.990 193.045 105.055 193.085 ;
        RECT 97.600 191.820 98.200 192.420 ;
        RECT 77.720 189.625 78.250 190.155 ;
        RECT 98.805 189.780 103.555 189.950 ;
        RECT 103.325 189.265 103.495 189.780 ;
        RECT 103.990 189.700 104.320 193.045 ;
        RECT 112.070 192.935 112.400 194.310 ;
        RECT 112.705 192.935 113.235 193.175 ;
        RECT 112.070 192.645 113.235 192.935 ;
        RECT 112.070 192.605 113.135 192.645 ;
        RECT 105.795 191.820 106.395 192.420 ;
        RECT 106.885 189.780 111.635 189.950 ;
        RECT 107.180 189.265 107.480 189.780 ;
        RECT 112.070 189.700 112.400 192.605 ;
        RECT 45.720 187.570 46.050 187.650 ;
        RECT 46.585 187.570 47.285 188.745 ;
        RECT 103.145 188.735 103.675 189.265 ;
        RECT 107.065 188.735 107.595 189.265 ;
        RECT 44.660 186.870 46.050 187.570 ;
        RECT 46.465 187.400 53.255 187.570 ;
        RECT 45.720 185.040 46.050 186.870 ;
        RECT 53.870 186.055 54.400 186.585 ;
        RECT 46.465 185.120 53.255 185.290 ;
        RECT 52.950 184.760 53.250 185.120 ;
        RECT 52.860 184.230 53.390 184.760 ;
        RECT 58.555 184.040 58.725 185.920 ;
        RECT 118.890 185.250 119.060 185.920 ;
        RECT 45.720 183.115 46.050 183.175 ;
        RECT 44.660 182.415 46.050 183.115 ;
        RECT 46.585 183.095 47.285 184.015 ;
        RECT 46.465 182.925 53.255 183.095 ;
        RECT 45.720 180.565 46.050 182.415 ;
        RECT 53.870 181.600 54.400 182.130 ;
        RECT 58.555 181.620 58.725 183.500 ;
        RECT 118.890 182.830 119.060 184.710 ;
        RECT 46.465 180.645 53.255 180.815 ;
        RECT 52.945 180.245 53.245 180.645 ;
        RECT 52.860 179.715 53.390 180.245 ;
        RECT 45.720 178.515 46.050 178.560 ;
        RECT 44.660 177.815 46.050 178.515 ;
        RECT 46.585 178.480 47.285 179.450 ;
        RECT 58.555 179.200 58.725 181.080 ;
        RECT 118.890 180.410 119.060 182.290 ;
        RECT 118.890 179.200 119.060 179.870 ;
        RECT 46.465 178.310 53.255 178.480 ;
        RECT 45.720 175.950 46.050 177.815 ;
        RECT 53.870 176.905 54.400 177.435 ;
        RECT 46.465 176.030 53.255 176.200 ;
        RECT 52.950 175.645 53.250 176.030 ;
        RECT 52.860 175.115 53.390 175.645 ;
        RECT 89.260 175.615 89.790 176.145 ;
        RECT 107.010 175.615 107.710 176.635 ;
        RECT 89.405 175.230 89.705 175.615 ;
        RECT 107.010 175.510 111.860 175.615 ;
        RECT 107.110 175.445 111.860 175.510 ;
        RECT 89.405 175.060 90.075 175.230 ;
        RECT 89.405 175.000 89.705 175.060 ;
        RECT 45.700 172.970 46.030 172.985 ;
        RECT 44.660 172.270 46.030 172.970 ;
        RECT 46.500 172.905 47.200 173.880 ;
        RECT 87.905 173.610 88.795 174.500 ;
        RECT 90.550 174.255 90.880 175.310 ;
        RECT 112.295 174.955 112.625 175.695 ;
        RECT 112.295 174.255 113.740 174.955 ;
        RECT 90.550 173.555 91.815 174.255 ;
        RECT 46.445 172.735 53.235 172.905 ;
        RECT 89.405 172.780 90.075 172.950 ;
        RECT 45.700 170.375 46.030 172.270 ;
        RECT 89.405 172.175 89.705 172.780 ;
        RECT 90.550 172.700 90.880 173.555 ;
        RECT 105.765 172.755 106.365 173.355 ;
        RECT 53.845 171.195 54.375 171.725 ;
        RECT 89.285 171.645 89.815 172.175 ;
        RECT 107.210 171.335 107.910 171.345 ;
        RECT 107.110 171.165 111.860 171.335 ;
        RECT 46.445 170.455 53.235 170.625 ;
        RECT 45.700 168.330 46.030 168.470 ;
        RECT 46.500 168.390 47.200 169.430 ;
        RECT 52.515 169.420 53.215 170.455 ;
        RECT 107.210 170.220 107.910 171.165 ;
        RECT 112.295 171.085 112.625 174.255 ;
        RECT 107.010 168.505 107.710 169.465 ;
        RECT 107.010 168.415 111.860 168.505 ;
        RECT 44.725 167.630 46.030 168.330 ;
        RECT 46.445 168.220 53.235 168.390 ;
        RECT 107.110 168.335 111.860 168.415 ;
        RECT 112.295 168.400 112.625 168.585 ;
        RECT 45.700 165.860 46.030 167.630 ;
        RECT 112.295 167.700 113.650 168.400 ;
        RECT 53.875 166.885 54.405 167.415 ;
        RECT 46.445 165.940 53.235 166.110 ;
        RECT 52.515 164.880 53.215 165.940 ;
        RECT 89.275 165.555 89.805 166.085 ;
        RECT 94.000 165.585 94.530 166.115 ;
        RECT 105.765 165.965 106.365 166.565 ;
        RECT 89.410 165.230 89.710 165.555 ;
        RECT 89.400 165.060 90.070 165.230 ;
        RECT 89.410 164.990 89.710 165.060 ;
        RECT 45.700 163.865 46.030 163.880 ;
        RECT 44.660 163.165 46.030 163.865 ;
        RECT 46.500 163.800 47.200 164.855 ;
        RECT 46.445 163.630 53.235 163.800 ;
        RECT 87.995 163.650 88.885 164.540 ;
        RECT 90.545 164.300 90.875 165.310 ;
        RECT 45.700 161.270 46.030 163.165 ;
        RECT 90.545 163.600 91.880 164.300 ;
        RECT 107.110 164.055 111.860 164.225 ;
        RECT 53.855 162.285 54.385 162.815 ;
        RECT 89.400 162.780 90.070 162.950 ;
        RECT 89.410 162.185 89.710 162.780 ;
        RECT 90.545 162.700 90.875 163.600 ;
        RECT 107.210 163.080 107.910 164.055 ;
        RECT 112.295 163.975 112.625 167.700 ;
        RECT 89.285 161.655 89.815 162.185 ;
        RECT 46.445 161.350 53.235 161.520 ;
        RECT 52.495 160.130 53.195 161.350 ;
        RECT 45.915 156.380 46.085 158.260 ;
        RECT 110.920 157.590 111.090 158.260 ;
        RECT 45.915 153.960 46.085 155.840 ;
        RECT 110.920 155.170 111.090 157.050 ;
        RECT 45.915 151.540 46.085 153.420 ;
        RECT 110.920 152.750 111.090 154.630 ;
        RECT 45.915 149.120 46.085 151.000 ;
        RECT 110.920 150.330 111.090 152.210 ;
        RECT 45.915 146.700 46.085 148.580 ;
        RECT 110.920 147.910 111.090 149.790 ;
        RECT 45.915 144.280 46.085 146.160 ;
        RECT 110.920 145.490 111.090 147.370 ;
        RECT 45.915 141.860 46.085 143.740 ;
        RECT 110.920 143.070 111.090 144.950 ;
        RECT 45.915 139.440 46.085 141.320 ;
        RECT 110.920 140.650 111.090 142.530 ;
        RECT 110.920 139.440 111.090 140.110 ;
        RECT 44.235 107.735 44.765 107.905 ;
        RECT 53.220 107.745 53.750 107.915 ;
        RECT 63.455 107.745 63.985 107.915 ;
        RECT 43.600 105.890 43.930 107.135 ;
        RECT 44.410 107.055 44.580 107.735 ;
        RECT 53.395 107.110 53.565 107.745 ;
        RECT 44.365 106.885 49.115 107.055 ;
        RECT 53.380 106.940 58.130 107.110 ;
        RECT 44.410 106.880 44.580 106.885 ;
        RECT 42.245 104.890 43.930 105.890 ;
        RECT 58.565 105.315 58.895 107.190 ;
        RECT 63.630 107.110 63.800 107.745 ;
        RECT 63.530 106.940 68.280 107.110 ;
        RECT 68.715 105.355 69.045 107.190 ;
        RECT 76.845 107.065 77.545 108.495 ;
        RECT 72.810 106.895 77.560 107.065 ;
        RECT 76.845 106.885 77.545 106.895 ;
        RECT 43.600 102.525 43.930 104.890 ;
        RECT 49.775 104.750 50.305 105.280 ;
        RECT 58.565 105.245 59.940 105.315 ;
        RECT 68.715 105.245 70.150 105.355 ;
        RECT 58.565 105.075 60.225 105.245 ;
        RECT 68.715 105.075 70.250 105.245 ;
        RECT 58.565 104.985 59.940 105.075 ;
        RECT 68.715 105.025 70.150 105.075 ;
        RECT 52.215 102.785 52.745 103.315 ;
        RECT 44.365 102.605 49.115 102.775 ;
        RECT 53.380 102.660 58.130 102.830 ;
        RECT 44.435 102.155 44.605 102.605 ;
        RECT 53.420 102.190 53.590 102.660 ;
        RECT 58.565 102.580 58.895 104.985 ;
        RECT 62.375 102.755 62.905 103.285 ;
        RECT 63.530 102.660 68.280 102.830 ;
        RECT 43.975 101.155 44.975 102.155 ;
        RECT 52.960 101.190 53.960 102.190 ;
        RECT 63.915 102.130 64.085 102.660 ;
        RECT 68.715 102.580 69.045 105.025 ;
        RECT 71.575 104.545 72.105 105.075 ;
        RECT 72.810 102.615 77.560 102.785 ;
        RECT 63.455 101.130 64.455 102.130 ;
        RECT 72.830 102.110 73.000 102.615 ;
        RECT 72.425 101.220 73.315 102.110 ;
        RECT 77.995 101.575 78.325 107.145 ;
        RECT 81.150 103.250 81.320 103.920 ;
        RECT 77.710 101.530 78.325 101.575 ;
        RECT 77.610 101.360 78.325 101.530 ;
        RECT 77.710 101.245 78.325 101.360 ;
        RECT 81.150 100.830 81.320 102.710 ;
        RECT 121.985 102.040 122.155 103.920 ;
        RECT 44.235 98.885 44.765 99.055 ;
        RECT 43.600 96.095 43.930 97.320 ;
        RECT 44.410 97.240 44.580 98.885 ;
        RECT 53.220 97.785 53.750 97.955 ;
        RECT 63.455 97.805 63.985 97.975 ;
        RECT 44.365 97.070 49.115 97.240 ;
        RECT 53.395 97.215 53.565 97.785 ;
        RECT 53.380 97.045 58.130 97.215 ;
        RECT 42.245 95.095 43.930 96.095 ;
        RECT 43.600 92.710 43.930 95.095 ;
        RECT 49.795 94.640 50.325 95.170 ;
        RECT 58.565 94.925 58.895 97.295 ;
        RECT 63.630 97.235 63.800 97.805 ;
        RECT 62.375 96.560 62.905 97.090 ;
        RECT 63.530 97.065 68.280 97.235 ;
        RECT 68.715 95.030 69.045 97.315 ;
        RECT 76.845 97.175 77.545 98.590 ;
        RECT 81.150 98.410 81.320 100.290 ;
        RECT 121.985 99.620 122.155 101.500 ;
        RECT 121.985 98.410 122.155 99.080 ;
        RECT 72.810 97.005 77.560 97.175 ;
        RECT 76.845 96.980 77.545 97.005 ;
        RECT 58.565 94.895 59.985 94.925 ;
        RECT 68.715 94.895 70.150 95.030 ;
        RECT 58.565 94.725 60.225 94.895 ;
        RECT 68.715 94.725 70.250 94.895 ;
        RECT 58.565 94.595 59.985 94.725 ;
        RECT 68.715 94.700 70.150 94.725 ;
        RECT 44.365 92.790 49.115 92.960 ;
        RECT 52.215 92.855 52.745 93.385 ;
        RECT 44.435 92.245 44.605 92.790 ;
        RECT 53.380 92.765 58.130 92.935 ;
        RECT 53.420 92.280 53.590 92.765 ;
        RECT 58.565 92.685 58.895 94.595 ;
        RECT 63.530 92.785 68.280 92.955 ;
        RECT 43.975 91.245 44.975 92.245 ;
        RECT 52.960 91.280 53.960 92.280 ;
        RECT 63.915 92.235 64.085 92.785 ;
        RECT 68.715 92.705 69.045 94.700 ;
        RECT 71.595 94.580 72.125 95.110 ;
        RECT 72.810 92.725 77.560 92.895 ;
        RECT 63.455 91.235 64.455 92.235 ;
        RECT 72.830 92.210 73.000 92.725 ;
        RECT 72.425 91.320 73.315 92.210 ;
        RECT 77.995 92.060 78.325 97.255 ;
        RECT 91.440 94.520 91.970 95.050 ;
        RECT 94.645 94.455 95.645 95.455 ;
        RECT 110.475 95.115 111.005 95.645 ;
        RECT 96.335 94.675 96.865 94.845 ;
        RECT 92.740 92.755 93.740 93.730 ;
        RECT 94.405 93.570 94.935 93.595 ;
        RECT 94.405 93.425 95.020 93.570 ;
        RECT 94.775 93.400 95.020 93.425 ;
        RECT 92.740 92.730 94.580 92.755 ;
        RECT 93.315 92.585 94.580 92.730 ;
        RECT 77.710 92.010 78.325 92.060 ;
        RECT 77.610 91.840 78.325 92.010 ;
        RECT 77.710 91.730 78.325 91.840 ;
        RECT 91.710 91.165 92.710 92.165 ;
        RECT 94.410 92.095 94.580 92.585 ;
        RECT 94.850 92.510 95.020 93.400 ;
        RECT 95.370 93.130 95.540 94.455 ;
        RECT 96.515 93.770 96.685 94.675 ;
        RECT 112.975 94.455 113.975 95.455 ;
        RECT 114.665 94.675 115.195 94.845 ;
        RECT 96.210 93.600 100.960 93.770 ;
        RECT 96.210 93.130 100.960 93.140 ;
        RECT 95.370 92.970 100.960 93.130 ;
        RECT 95.370 92.960 96.340 92.970 ;
        RECT 101.395 92.605 101.725 93.850 ;
        RECT 102.775 92.605 103.775 93.045 ;
        RECT 111.070 92.755 112.070 93.730 ;
        RECT 112.735 93.570 113.265 93.595 ;
        RECT 112.735 93.425 113.350 93.570 ;
        RECT 113.105 93.400 113.350 93.425 ;
        RECT 111.070 92.730 112.910 92.755 ;
        RECT 94.850 92.340 100.960 92.510 ;
        RECT 101.395 92.275 103.775 92.605 ;
        RECT 111.645 92.585 112.910 92.730 ;
        RECT 94.410 91.925 95.910 92.095 ;
        RECT 93.355 91.755 93.970 91.925 ;
        RECT 93.800 91.690 93.970 91.755 ;
        RECT 95.740 91.880 95.910 91.925 ;
        RECT 95.740 91.710 100.960 91.880 ;
        RECT 93.800 91.520 95.450 91.690 ;
        RECT 95.280 91.450 95.450 91.520 ;
        RECT 95.280 91.280 95.925 91.450 ;
        RECT 92.540 91.060 92.710 91.165 ;
        RECT 95.755 91.250 95.925 91.280 ;
        RECT 95.755 91.080 100.960 91.250 ;
        RECT 92.540 90.890 95.345 91.060 ;
        RECT 89.360 89.660 90.360 90.660 ;
        RECT 95.175 90.620 95.345 90.890 ;
        RECT 91.600 90.410 94.985 90.580 ;
        RECT 95.175 90.450 100.960 90.620 ;
        RECT 91.600 90.345 91.770 90.410 ;
        RECT 91.240 90.175 91.770 90.345 ;
        RECT 92.395 89.885 94.260 90.055 ;
        RECT 88.040 89.445 88.570 89.530 ;
        RECT 88.040 89.275 88.830 89.445 ;
        RECT 88.660 88.875 88.830 89.275 ;
        RECT 90.010 89.335 90.180 89.660 ;
        RECT 92.395 89.335 92.565 89.885 ;
        RECT 90.010 89.165 92.565 89.335 ;
        RECT 94.090 89.360 94.260 89.885 ;
        RECT 94.815 89.990 94.985 90.410 ;
        RECT 94.815 89.820 100.960 89.990 ;
        RECT 94.090 89.190 100.960 89.360 ;
        RECT 89.650 88.875 91.925 88.900 ;
        RECT 53.220 88.015 53.750 88.185 ;
        RECT 63.455 88.140 63.985 88.310 ;
        RECT 44.235 87.665 44.765 87.835 ;
        RECT 43.600 86.735 43.930 87.160 ;
        RECT 44.410 87.080 44.580 87.665 ;
        RECT 53.405 87.170 53.575 88.015 ;
        RECT 63.640 87.295 63.810 88.140 ;
        RECT 44.365 86.910 49.115 87.080 ;
        RECT 53.380 87.000 58.130 87.170 ;
        RECT 42.245 85.735 43.930 86.735 ;
        RECT 43.600 82.550 43.930 85.735 ;
        RECT 49.775 84.565 50.305 85.095 ;
        RECT 58.565 84.940 58.895 87.250 ;
        RECT 63.530 87.125 68.280 87.295 ;
        RECT 62.375 86.555 62.905 87.085 ;
        RECT 68.715 85.090 69.045 87.375 ;
        RECT 76.795 87.340 77.495 88.780 ;
        RECT 88.660 88.730 91.925 88.875 ;
        RECT 88.660 88.705 89.820 88.730 ;
        RECT 91.755 88.560 100.960 88.730 ;
        RECT 86.145 88.100 87.145 88.500 ;
        RECT 86.145 87.930 100.960 88.100 ;
        RECT 86.145 87.500 87.145 87.930 ;
        RECT 96.210 87.440 100.960 87.470 ;
        RECT 72.765 87.170 77.515 87.340 ;
        RECT 68.715 85.035 70.150 85.090 ;
        RECT 58.565 84.875 60.030 84.940 ;
        RECT 58.565 84.705 60.225 84.875 ;
        RECT 68.715 84.865 70.250 85.035 ;
        RECT 68.715 84.760 70.150 84.865 ;
        RECT 71.535 84.820 72.065 85.350 ;
        RECT 58.565 84.610 60.030 84.705 ;
        RECT 52.215 82.805 52.745 83.335 ;
        RECT 44.365 82.630 49.115 82.800 ;
        RECT 53.380 82.720 58.130 82.890 ;
        RECT 44.435 82.090 44.605 82.630 ;
        RECT 53.420 82.265 53.590 82.720 ;
        RECT 58.565 82.640 58.895 84.610 ;
        RECT 63.530 82.845 68.280 83.015 ;
        RECT 63.915 82.380 64.085 82.845 ;
        RECT 68.715 82.765 69.045 84.760 ;
        RECT 72.765 82.890 77.515 83.060 ;
        RECT 72.770 82.530 72.940 82.890 ;
        RECT 43.975 81.090 44.975 82.090 ;
        RECT 52.960 81.265 53.960 82.265 ;
        RECT 63.455 81.380 64.455 82.380 ;
        RECT 72.500 81.530 73.500 82.530 ;
        RECT 77.950 81.655 78.280 87.420 ;
        RECT 94.670 87.300 100.960 87.440 ;
        RECT 94.670 87.270 96.425 87.300 ;
        RECT 94.670 87.170 94.840 87.270 ;
        RECT 88.040 87.000 94.840 87.170 ;
        RECT 95.235 86.840 96.375 86.855 ;
        RECT 95.235 86.685 100.960 86.840 ;
        RECT 95.235 86.635 95.405 86.685 ;
        RECT 96.210 86.670 100.960 86.685 ;
        RECT 89.095 86.465 95.405 86.635 ;
        RECT 89.095 86.120 89.265 86.465 ;
        RECT 96.210 86.190 100.960 86.210 ;
        RECT 95.695 86.150 100.960 86.190 ;
        RECT 88.680 85.120 89.680 86.120 ;
        RECT 90.820 86.040 100.960 86.150 ;
        RECT 90.820 86.020 96.365 86.040 ;
        RECT 90.820 85.980 95.865 86.020 ;
        RECT 90.820 85.705 90.990 85.980 ;
        RECT 90.375 85.535 90.990 85.705 ;
        RECT 91.475 85.410 100.960 85.580 ;
        RECT 91.475 84.695 91.645 85.410 ;
        RECT 92.940 84.780 100.960 84.950 ;
        RECT 90.755 83.695 91.755 84.695 ;
        RECT 92.940 84.185 93.110 84.780 ;
        RECT 92.480 84.015 93.110 84.185 ;
        RECT 92.660 83.975 93.110 84.015 ;
        RECT 93.650 84.150 100.960 84.320 ;
        RECT 93.650 83.280 93.820 84.150 ;
        RECT 91.630 83.110 93.820 83.280 ;
        RECT 94.260 83.520 100.960 83.690 ;
        RECT 91.630 82.750 91.800 83.110 ;
        RECT 90.755 82.165 91.800 82.750 ;
        RECT 94.260 82.430 94.430 83.520 ;
        RECT 92.865 82.360 94.430 82.430 ;
        RECT 92.685 82.260 94.430 82.360 ;
        RECT 94.880 82.890 100.960 83.060 ;
        RECT 92.685 82.190 93.215 82.260 ;
        RECT 90.755 81.750 91.755 82.165 ;
        RECT 94.880 81.875 95.050 82.890 ;
        RECT 77.575 81.490 78.280 81.655 ;
        RECT 93.820 81.705 95.050 81.875 ;
        RECT 95.370 82.260 100.960 82.430 ;
        RECT 77.575 81.485 78.105 81.490 ;
        RECT 93.820 81.210 93.990 81.705 ;
        RECT 93.025 80.210 94.025 81.210 ;
        RECT 95.370 80.935 95.540 82.260 ;
        RECT 96.210 81.630 100.960 81.800 ;
        RECT 96.595 81.210 96.765 81.630 ;
        RECT 101.395 81.550 101.725 92.275 ;
        RECT 102.775 92.045 103.775 92.275 ;
        RECT 110.040 91.165 111.040 92.165 ;
        RECT 112.740 92.095 112.910 92.585 ;
        RECT 113.180 92.510 113.350 93.400 ;
        RECT 113.700 93.130 113.870 94.455 ;
        RECT 114.845 93.770 115.015 94.675 ;
        RECT 114.555 93.600 119.305 93.770 ;
        RECT 114.555 93.130 119.305 93.140 ;
        RECT 113.700 92.970 119.305 93.130 ;
        RECT 113.700 92.960 114.670 92.970 ;
        RECT 113.180 92.340 119.305 92.510 ;
        RECT 112.740 91.925 114.240 92.095 ;
        RECT 111.685 91.755 112.300 91.925 ;
        RECT 112.130 91.690 112.300 91.755 ;
        RECT 114.070 91.880 114.240 91.925 ;
        RECT 114.070 91.710 119.305 91.880 ;
        RECT 112.130 91.520 113.780 91.690 ;
        RECT 113.610 91.450 113.780 91.520 ;
        RECT 113.610 91.280 114.255 91.450 ;
        RECT 110.870 91.060 111.040 91.165 ;
        RECT 114.085 91.250 114.255 91.280 ;
        RECT 114.085 91.080 119.305 91.250 ;
        RECT 110.870 90.890 113.675 91.060 ;
        RECT 107.690 89.660 108.690 90.660 ;
        RECT 113.505 90.620 113.675 90.890 ;
        RECT 109.930 90.410 113.315 90.580 ;
        RECT 113.505 90.450 119.305 90.620 ;
        RECT 109.930 90.345 110.100 90.410 ;
        RECT 109.570 90.175 110.100 90.345 ;
        RECT 110.725 89.885 112.590 90.055 ;
        RECT 106.370 89.445 106.900 89.530 ;
        RECT 106.370 89.275 107.160 89.445 ;
        RECT 106.990 88.875 107.160 89.275 ;
        RECT 108.340 89.335 108.510 89.660 ;
        RECT 110.725 89.335 110.895 89.885 ;
        RECT 108.340 89.165 110.895 89.335 ;
        RECT 112.420 89.360 112.590 89.885 ;
        RECT 113.145 89.990 113.315 90.410 ;
        RECT 113.145 89.820 119.305 89.990 ;
        RECT 112.420 89.190 119.305 89.360 ;
        RECT 107.980 88.875 110.255 88.900 ;
        RECT 106.990 88.730 110.255 88.875 ;
        RECT 106.990 88.705 108.150 88.730 ;
        RECT 110.085 88.560 119.305 88.730 ;
        RECT 104.475 88.100 105.475 88.520 ;
        RECT 119.740 88.475 120.070 93.850 ;
        RECT 104.475 87.930 119.305 88.100 ;
        RECT 104.475 87.520 105.475 87.930 ;
        RECT 119.740 87.775 121.185 88.475 ;
        RECT 114.555 87.440 119.305 87.470 ;
        RECT 113.000 87.300 119.305 87.440 ;
        RECT 113.000 87.270 114.755 87.300 ;
        RECT 113.000 87.170 113.170 87.270 ;
        RECT 106.370 87.000 113.170 87.170 ;
        RECT 113.565 86.840 114.705 86.855 ;
        RECT 113.565 86.685 119.305 86.840 ;
        RECT 113.565 86.635 113.735 86.685 ;
        RECT 114.555 86.670 119.305 86.685 ;
        RECT 107.425 86.465 113.735 86.635 ;
        RECT 107.425 86.120 107.595 86.465 ;
        RECT 114.555 86.190 119.305 86.210 ;
        RECT 114.025 86.150 119.305 86.190 ;
        RECT 107.010 85.120 108.010 86.120 ;
        RECT 109.150 86.040 119.305 86.150 ;
        RECT 109.150 86.020 114.695 86.040 ;
        RECT 109.150 85.980 114.195 86.020 ;
        RECT 109.150 85.705 109.320 85.980 ;
        RECT 108.705 85.535 109.320 85.705 ;
        RECT 109.805 85.410 119.305 85.580 ;
        RECT 109.805 84.695 109.975 85.410 ;
        RECT 111.270 84.780 119.305 84.950 ;
        RECT 109.085 83.695 110.085 84.695 ;
        RECT 111.270 84.185 111.440 84.780 ;
        RECT 110.810 84.015 111.440 84.185 ;
        RECT 110.990 83.975 111.440 84.015 ;
        RECT 111.980 84.150 119.305 84.320 ;
        RECT 111.980 83.280 112.150 84.150 ;
        RECT 109.960 83.110 112.150 83.280 ;
        RECT 112.590 83.520 119.305 83.690 ;
        RECT 109.960 82.750 110.130 83.110 ;
        RECT 109.085 82.165 110.130 82.750 ;
        RECT 112.590 82.430 112.760 83.520 ;
        RECT 111.195 82.360 112.760 82.430 ;
        RECT 111.015 82.260 112.760 82.360 ;
        RECT 113.210 82.890 119.305 83.060 ;
        RECT 111.015 82.190 111.545 82.260 ;
        RECT 109.085 81.750 110.085 82.165 ;
        RECT 113.210 81.875 113.380 82.890 ;
        RECT 112.150 81.705 113.380 81.875 ;
        RECT 113.700 82.260 119.305 82.430 ;
        RECT 112.150 81.210 112.320 81.705 ;
        RECT 94.945 80.900 95.540 80.935 ;
        RECT 94.765 80.765 95.540 80.900 ;
        RECT 94.765 80.730 95.295 80.765 ;
        RECT 96.180 80.210 97.180 81.210 ;
        RECT 111.355 80.210 112.355 81.210 ;
        RECT 113.700 80.935 113.870 82.260 ;
        RECT 114.555 81.630 119.305 81.800 ;
        RECT 114.925 81.210 115.095 81.630 ;
        RECT 119.740 81.550 120.070 87.775 ;
        RECT 113.275 80.900 113.870 80.935 ;
        RECT 113.095 80.765 113.870 80.900 ;
        RECT 113.095 80.730 113.625 80.765 ;
        RECT 114.510 80.210 115.510 81.210 ;
        RECT 44.235 78.590 44.765 78.760 ;
        RECT 43.600 76.165 43.930 78.095 ;
        RECT 44.410 78.015 44.580 78.590 ;
        RECT 53.220 78.580 53.750 78.750 ;
        RECT 63.455 78.625 63.985 78.795 ;
        RECT 44.365 77.845 49.115 78.015 ;
        RECT 53.395 77.970 53.565 78.580 ;
        RECT 52.215 77.385 52.745 77.915 ;
        RECT 53.380 77.800 58.130 77.970 ;
        RECT 41.875 75.165 43.930 76.165 ;
        RECT 58.565 75.990 58.895 78.050 ;
        RECT 63.630 77.875 63.800 78.625 ;
        RECT 77.045 78.480 77.575 78.485 ;
        RECT 76.865 78.315 77.575 78.480 ;
        RECT 62.375 77.290 62.905 77.820 ;
        RECT 63.530 77.705 68.280 77.875 ;
        RECT 58.565 75.940 59.995 75.990 ;
        RECT 49.795 75.365 50.325 75.895 ;
        RECT 58.565 75.770 60.225 75.940 ;
        RECT 58.565 75.660 59.995 75.770 ;
        RECT 68.715 75.760 69.045 77.955 ;
        RECT 76.865 77.780 77.565 78.315 ;
        RECT 72.810 77.610 77.565 77.780 ;
        RECT 76.865 77.595 77.565 77.610 ;
        RECT 68.715 75.710 69.925 75.760 ;
        RECT 43.600 73.485 43.930 75.165 ;
        RECT 44.365 73.565 49.115 73.735 ;
        RECT 44.435 73.085 44.605 73.565 ;
        RECT 53.380 73.520 58.130 73.690 ;
        RECT 43.975 72.085 44.975 73.085 ;
        RECT 53.420 73.060 53.590 73.520 ;
        RECT 58.565 73.440 58.895 75.660 ;
        RECT 68.715 75.540 70.250 75.710 ;
        RECT 68.715 75.430 69.925 75.540 ;
        RECT 63.530 73.425 68.280 73.595 ;
        RECT 63.915 73.205 64.085 73.425 ;
        RECT 68.715 73.345 69.045 75.430 ;
        RECT 71.555 75.120 72.085 75.650 ;
        RECT 72.820 73.500 72.990 73.520 ;
        RECT 72.810 73.330 77.560 73.500 ;
        RECT 52.960 72.060 53.960 73.060 ;
        RECT 63.455 72.205 64.455 73.205 ;
        RECT 72.820 72.905 72.990 73.330 ;
        RECT 72.095 71.905 73.095 72.905 ;
        RECT 77.995 72.215 78.325 77.860 ;
        RECT 91.130 76.135 91.660 76.665 ;
        RECT 94.405 76.165 95.405 77.165 ;
        RECT 96.045 76.385 96.575 76.555 ;
        RECT 92.450 74.465 93.450 75.440 ;
        RECT 94.115 75.280 94.645 75.305 ;
        RECT 94.115 75.135 94.730 75.280 ;
        RECT 94.485 75.110 94.730 75.135 ;
        RECT 92.450 74.440 94.290 74.465 ;
        RECT 93.025 74.295 94.290 74.440 ;
        RECT 91.420 72.875 92.420 73.875 ;
        RECT 94.120 73.805 94.290 74.295 ;
        RECT 94.560 74.220 94.730 75.110 ;
        RECT 95.080 74.840 95.250 76.165 ;
        RECT 96.225 75.480 96.395 76.385 ;
        RECT 109.780 75.760 110.310 76.290 ;
        RECT 113.005 75.920 114.005 76.920 ;
        RECT 114.695 76.140 115.225 76.310 ;
        RECT 95.905 75.310 100.655 75.480 ;
        RECT 95.905 74.840 100.655 74.850 ;
        RECT 95.080 74.680 100.655 74.840 ;
        RECT 95.080 74.670 96.050 74.680 ;
        RECT 94.560 74.050 100.655 74.220 ;
        RECT 94.120 73.635 95.620 73.805 ;
        RECT 93.065 73.465 93.680 73.635 ;
        RECT 93.510 73.400 93.680 73.465 ;
        RECT 95.450 73.590 95.620 73.635 ;
        RECT 95.450 73.420 100.655 73.590 ;
        RECT 93.510 73.230 95.160 73.400 ;
        RECT 94.990 73.160 95.160 73.230 ;
        RECT 94.990 72.990 95.635 73.160 ;
        RECT 92.250 72.770 92.420 72.875 ;
        RECT 95.465 72.960 95.635 72.990 ;
        RECT 95.465 72.790 100.655 72.960 ;
        RECT 92.250 72.600 95.055 72.770 ;
        RECT 77.705 71.885 78.325 72.215 ;
        RECT 89.070 71.370 90.070 72.370 ;
        RECT 94.885 72.330 95.055 72.600 ;
        RECT 91.310 72.120 94.695 72.290 ;
        RECT 94.885 72.160 100.655 72.330 ;
        RECT 91.310 72.055 91.480 72.120 ;
        RECT 90.950 71.885 91.480 72.055 ;
        RECT 92.105 71.595 93.970 71.765 ;
        RECT 87.750 71.155 88.280 71.240 ;
        RECT 87.750 70.985 88.540 71.155 ;
        RECT 49.285 70.755 50.350 70.850 ;
        RECT 49.285 70.585 50.450 70.755 ;
        RECT 88.370 70.585 88.540 70.985 ;
        RECT 89.720 71.045 89.890 71.370 ;
        RECT 92.105 71.045 92.275 71.595 ;
        RECT 89.720 70.875 92.275 71.045 ;
        RECT 93.800 71.070 93.970 71.595 ;
        RECT 94.525 71.700 94.695 72.120 ;
        RECT 94.525 71.530 100.655 71.700 ;
        RECT 93.800 70.900 100.655 71.070 ;
        RECT 89.360 70.585 91.635 70.610 ;
        RECT 49.285 70.520 50.350 70.585 ;
        RECT 49.285 66.270 49.615 70.520 ;
        RECT 50.050 69.800 50.220 70.520 ;
        RECT 88.370 70.440 91.635 70.585 ;
        RECT 88.370 70.415 89.530 70.440 ;
        RECT 91.465 70.270 100.655 70.440 ;
        RECT 85.855 69.810 86.855 70.230 ;
        RECT 50.040 69.630 55.810 69.800 ;
        RECT 85.855 69.640 100.655 69.810 ;
        RECT 85.855 69.230 86.855 69.640 ;
        RECT 95.905 69.150 100.655 69.180 ;
        RECT 94.380 69.010 100.655 69.150 ;
        RECT 94.380 68.980 96.135 69.010 ;
        RECT 94.380 68.880 94.550 68.980 ;
        RECT 87.750 68.710 94.550 68.880 ;
        RECT 94.945 68.550 96.085 68.565 ;
        RECT 73.840 68.255 74.370 68.430 ;
        RECT 94.945 68.395 100.655 68.550 ;
        RECT 94.945 68.345 95.115 68.395 ;
        RECT 95.905 68.380 100.655 68.395 ;
        RECT 73.840 68.085 81.850 68.255 ;
        RECT 73.840 67.900 74.370 68.085 ;
        RECT 62.095 67.785 62.825 67.790 ;
        RECT 61.915 67.775 62.825 67.785 ;
        RECT 56.450 67.110 56.980 67.640 ;
        RECT 61.915 67.620 69.495 67.775 ;
        RECT 61.915 67.615 62.445 67.620 ;
        RECT 62.705 67.605 69.495 67.620 ;
        RECT 59.765 66.695 69.495 66.865 ;
        RECT 50.040 66.500 55.810 66.520 ;
        RECT 50.030 66.350 55.810 66.500 ;
        RECT 50.030 65.885 50.200 66.350 ;
        RECT 49.570 64.885 50.570 65.885 ;
        RECT 59.765 65.045 59.935 66.695 ;
        RECT 62.095 65.965 62.955 65.970 ;
        RECT 61.915 65.955 62.955 65.965 ;
        RECT 61.915 65.800 69.495 65.955 ;
        RECT 61.915 65.795 62.445 65.800 ;
        RECT 62.705 65.785 69.495 65.800 ;
        RECT 59.765 64.875 69.495 65.045 ;
        RECT 49.285 64.215 50.350 64.245 ;
        RECT 49.285 64.045 50.450 64.215 ;
        RECT 49.285 63.915 50.350 64.045 ;
        RECT 49.285 59.580 49.615 63.915 ;
        RECT 50.040 63.110 50.210 63.915 ;
        RECT 59.765 63.225 59.935 64.875 ;
        RECT 62.095 64.145 62.935 64.150 ;
        RECT 61.915 64.135 62.935 64.145 ;
        RECT 61.915 63.980 69.495 64.135 ;
        RECT 61.915 63.975 62.445 63.980 ;
        RECT 62.705 63.965 69.495 63.980 ;
        RECT 50.040 62.940 55.810 63.110 ;
        RECT 59.765 63.055 69.495 63.225 ;
        RECT 56.470 61.775 57.000 62.305 ;
        RECT 59.765 61.405 59.935 63.055 ;
        RECT 61.925 62.315 62.825 62.330 ;
        RECT 61.925 62.160 69.495 62.315 ;
        RECT 62.705 62.145 69.495 62.160 ;
        RECT 59.765 61.235 69.495 61.405 ;
        RECT 50.040 59.810 55.810 59.830 ;
        RECT 50.030 59.660 55.810 59.810 ;
        RECT 50.030 59.195 50.200 59.660 ;
        RECT 59.765 59.585 59.935 61.235 ;
        RECT 61.925 60.495 62.455 60.505 ;
        RECT 61.925 60.335 69.495 60.495 ;
        RECT 62.105 60.325 69.495 60.335 ;
        RECT 59.765 59.415 69.495 59.585 ;
        RECT 49.570 58.195 50.570 59.195 ;
        RECT 59.765 57.765 59.935 59.415 ;
        RECT 62.105 58.680 62.970 58.690 ;
        RECT 61.925 58.675 62.970 58.680 ;
        RECT 61.925 58.520 69.495 58.675 ;
        RECT 61.925 58.510 62.455 58.520 ;
        RECT 62.705 58.505 69.495 58.520 ;
        RECT 59.765 57.595 69.495 57.765 ;
        RECT 49.285 57.520 50.350 57.590 ;
        RECT 49.285 57.350 50.450 57.520 ;
        RECT 49.285 57.260 50.350 57.350 ;
        RECT 49.285 52.890 49.615 57.260 ;
        RECT 50.045 56.420 50.215 57.260 ;
        RECT 59.765 56.755 59.935 57.595 ;
        RECT 61.915 56.855 62.960 56.870 ;
        RECT 60.335 56.755 60.605 56.840 ;
        RECT 59.765 56.585 60.605 56.755 ;
        RECT 61.915 56.700 69.495 56.855 ;
        RECT 62.705 56.685 69.495 56.700 ;
        RECT 50.040 56.250 55.810 56.420 ;
        RECT 59.765 55.945 59.935 56.585 ;
        RECT 60.335 56.510 60.605 56.585 ;
        RECT 59.765 55.775 69.495 55.945 ;
        RECT 59.765 55.045 59.935 55.775 ;
        RECT 62.190 55.050 62.385 55.165 ;
        RECT 62.190 55.045 62.920 55.050 ;
        RECT 59.620 54.875 60.150 55.045 ;
        RECT 61.925 55.035 62.920 55.045 ;
        RECT 61.925 54.880 69.495 55.035 ;
        RECT 69.910 55.020 70.240 67.855 ;
        RECT 72.640 66.805 81.850 66.975 ;
        RECT 72.690 64.415 72.860 66.805 ;
        RECT 73.840 65.695 74.370 65.915 ;
        RECT 73.840 65.525 81.850 65.695 ;
        RECT 73.840 65.385 74.370 65.525 ;
        RECT 72.690 64.245 81.850 64.415 ;
        RECT 72.690 61.855 72.860 64.245 ;
        RECT 73.840 63.135 74.370 63.310 ;
        RECT 73.840 62.965 81.850 63.135 ;
        RECT 73.840 62.780 74.370 62.965 ;
        RECT 72.690 61.685 81.850 61.855 ;
        RECT 72.690 59.295 72.860 61.685 ;
        RECT 73.840 60.575 74.370 60.780 ;
        RECT 73.840 60.405 81.850 60.575 ;
        RECT 73.840 60.250 74.370 60.405 ;
        RECT 72.690 59.125 81.850 59.295 ;
        RECT 72.690 56.735 72.860 59.125 ;
        RECT 73.840 58.015 74.370 58.135 ;
        RECT 73.840 57.845 81.850 58.015 ;
        RECT 73.840 57.605 74.370 57.845 ;
        RECT 72.690 56.565 81.850 56.735 ;
        RECT 72.690 56.155 72.860 56.565 ;
        RECT 72.690 56.005 72.965 56.155 ;
        RECT 72.695 55.825 72.965 56.005 ;
        RECT 61.925 54.875 62.455 54.880 ;
        RECT 62.705 54.865 69.495 54.880 ;
        RECT 69.890 54.785 70.240 55.020 ;
        RECT 72.720 54.990 72.890 55.825 ;
        RECT 73.840 55.455 74.370 55.660 ;
        RECT 73.840 55.285 81.850 55.455 ;
        RECT 73.840 55.130 74.370 55.285 ;
        RECT 82.265 55.205 82.595 68.335 ;
        RECT 88.805 68.175 95.115 68.345 ;
        RECT 88.805 67.830 88.975 68.175 ;
        RECT 95.905 67.900 100.655 67.920 ;
        RECT 95.405 67.860 100.655 67.900 ;
        RECT 88.390 66.830 89.390 67.830 ;
        RECT 90.530 67.750 100.655 67.860 ;
        RECT 90.530 67.730 96.075 67.750 ;
        RECT 90.530 67.690 95.575 67.730 ;
        RECT 90.530 67.415 90.700 67.690 ;
        RECT 90.085 67.245 90.700 67.415 ;
        RECT 91.185 67.120 100.655 67.290 ;
        RECT 91.185 66.405 91.355 67.120 ;
        RECT 92.650 66.490 100.655 66.660 ;
        RECT 90.465 65.405 91.465 66.405 ;
        RECT 92.650 65.895 92.820 66.490 ;
        RECT 92.190 65.725 92.820 65.895 ;
        RECT 92.370 65.685 92.820 65.725 ;
        RECT 93.360 65.860 100.655 66.030 ;
        RECT 93.360 64.990 93.530 65.860 ;
        RECT 91.340 64.820 93.530 64.990 ;
        RECT 93.970 65.230 100.655 65.400 ;
        RECT 91.340 64.460 91.510 64.820 ;
        RECT 90.465 63.875 91.510 64.460 ;
        RECT 93.970 64.140 94.140 65.230 ;
        RECT 92.575 64.070 94.140 64.140 ;
        RECT 92.395 63.970 94.140 64.070 ;
        RECT 94.590 64.600 100.655 64.770 ;
        RECT 92.395 63.900 92.925 63.970 ;
        RECT 90.465 63.460 91.465 63.875 ;
        RECT 94.590 63.585 94.760 64.600 ;
        RECT 101.090 64.315 101.420 75.560 ;
        RECT 111.100 74.220 112.100 75.195 ;
        RECT 112.765 75.035 113.295 75.060 ;
        RECT 112.765 74.890 113.380 75.035 ;
        RECT 113.135 74.865 113.380 74.890 ;
        RECT 111.100 74.195 112.940 74.220 ;
        RECT 111.675 74.050 112.940 74.195 ;
        RECT 110.070 72.630 111.070 73.630 ;
        RECT 112.770 73.560 112.940 74.050 ;
        RECT 113.210 73.975 113.380 74.865 ;
        RECT 113.730 74.595 113.900 75.920 ;
        RECT 114.875 75.235 115.045 76.140 ;
        RECT 114.560 75.065 119.310 75.235 ;
        RECT 114.560 74.595 119.310 74.605 ;
        RECT 113.730 74.435 119.310 74.595 ;
        RECT 113.730 74.425 114.700 74.435 ;
        RECT 113.210 73.805 119.310 73.975 ;
        RECT 112.770 73.390 114.270 73.560 ;
        RECT 111.715 73.220 112.330 73.390 ;
        RECT 112.160 73.155 112.330 73.220 ;
        RECT 114.100 73.345 114.270 73.390 ;
        RECT 114.100 73.175 119.310 73.345 ;
        RECT 112.160 72.985 113.810 73.155 ;
        RECT 113.640 72.915 113.810 72.985 ;
        RECT 113.640 72.745 114.285 72.915 ;
        RECT 110.900 72.525 111.070 72.630 ;
        RECT 114.115 72.715 114.285 72.745 ;
        RECT 114.115 72.545 119.310 72.715 ;
        RECT 110.900 72.355 113.705 72.525 ;
        RECT 107.720 71.125 108.720 72.125 ;
        RECT 113.535 72.085 113.705 72.355 ;
        RECT 109.960 71.875 113.345 72.045 ;
        RECT 113.535 71.915 119.310 72.085 ;
        RECT 109.960 71.810 110.130 71.875 ;
        RECT 109.600 71.640 110.130 71.810 ;
        RECT 110.755 71.350 112.620 71.520 ;
        RECT 106.400 70.910 106.930 70.995 ;
        RECT 106.400 70.740 107.190 70.910 ;
        RECT 107.020 70.340 107.190 70.740 ;
        RECT 108.370 70.800 108.540 71.125 ;
        RECT 110.755 70.800 110.925 71.350 ;
        RECT 108.370 70.630 110.925 70.800 ;
        RECT 112.450 70.825 112.620 71.350 ;
        RECT 113.175 71.455 113.345 71.875 ;
        RECT 113.175 71.285 119.310 71.455 ;
        RECT 112.450 70.655 119.310 70.825 ;
        RECT 108.010 70.340 110.285 70.365 ;
        RECT 107.020 70.195 110.285 70.340 ;
        RECT 107.020 70.170 108.180 70.195 ;
        RECT 110.115 70.025 119.310 70.195 ;
        RECT 104.505 69.565 105.505 70.000 ;
        RECT 119.745 69.870 120.075 75.315 ;
        RECT 104.505 69.395 119.310 69.565 ;
        RECT 104.505 69.000 105.505 69.395 ;
        RECT 119.745 69.170 120.910 69.870 ;
        RECT 114.560 68.905 119.310 68.935 ;
        RECT 113.030 68.765 119.310 68.905 ;
        RECT 113.030 68.735 114.785 68.765 ;
        RECT 113.030 68.635 113.200 68.735 ;
        RECT 106.400 68.465 113.200 68.635 ;
        RECT 113.595 68.305 114.735 68.320 ;
        RECT 113.595 68.150 119.310 68.305 ;
        RECT 113.595 68.100 113.765 68.150 ;
        RECT 114.560 68.135 119.310 68.150 ;
        RECT 107.455 67.930 113.765 68.100 ;
        RECT 107.455 67.585 107.625 67.930 ;
        RECT 114.560 67.655 119.310 67.675 ;
        RECT 114.055 67.615 119.310 67.655 ;
        RECT 107.040 66.585 108.040 67.585 ;
        RECT 109.180 67.505 119.310 67.615 ;
        RECT 109.180 67.485 114.725 67.505 ;
        RECT 109.180 67.445 114.225 67.485 ;
        RECT 109.180 67.170 109.350 67.445 ;
        RECT 108.735 67.000 109.350 67.170 ;
        RECT 109.835 66.875 119.310 67.045 ;
        RECT 109.835 66.160 110.005 66.875 ;
        RECT 111.300 66.245 119.310 66.415 ;
        RECT 109.115 65.160 110.115 66.160 ;
        RECT 111.300 65.650 111.470 66.245 ;
        RECT 110.840 65.480 111.470 65.650 ;
        RECT 111.020 65.440 111.470 65.480 ;
        RECT 112.010 65.615 119.310 65.785 ;
        RECT 112.010 64.745 112.180 65.615 ;
        RECT 109.990 64.575 112.180 64.745 ;
        RECT 112.620 64.985 119.310 65.155 ;
        RECT 102.280 64.315 102.810 64.430 ;
        RECT 93.530 63.415 94.760 63.585 ;
        RECT 95.080 63.970 100.655 64.140 ;
        RECT 101.090 64.015 102.810 64.315 ;
        RECT 109.990 64.215 110.160 64.575 ;
        RECT 93.530 62.920 93.700 63.415 ;
        RECT 92.735 61.920 93.735 62.920 ;
        RECT 95.080 62.645 95.250 63.970 ;
        RECT 95.905 63.340 100.655 63.510 ;
        RECT 96.305 62.920 96.475 63.340 ;
        RECT 101.090 63.260 101.420 64.015 ;
        RECT 102.280 63.900 102.810 64.015 ;
        RECT 109.115 63.630 110.160 64.215 ;
        RECT 112.620 63.895 112.790 64.985 ;
        RECT 111.225 63.825 112.790 63.895 ;
        RECT 111.045 63.725 112.790 63.825 ;
        RECT 113.240 64.355 119.310 64.525 ;
        RECT 111.045 63.655 111.575 63.725 ;
        RECT 109.115 63.215 110.115 63.630 ;
        RECT 113.240 63.340 113.410 64.355 ;
        RECT 112.180 63.170 113.410 63.340 ;
        RECT 113.730 63.725 119.310 63.895 ;
        RECT 94.655 62.610 95.250 62.645 ;
        RECT 94.475 62.475 95.250 62.610 ;
        RECT 94.475 62.440 95.005 62.475 ;
        RECT 95.890 61.920 96.890 62.920 ;
        RECT 112.180 62.675 112.350 63.170 ;
        RECT 111.385 61.675 112.385 62.675 ;
        RECT 113.730 62.400 113.900 63.725 ;
        RECT 114.560 63.095 119.310 63.265 ;
        RECT 114.955 62.675 115.125 63.095 ;
        RECT 119.745 63.015 120.075 69.170 ;
        RECT 113.305 62.365 113.900 62.400 ;
        RECT 113.125 62.230 113.900 62.365 ;
        RECT 113.125 62.195 113.655 62.230 ;
        RECT 114.540 61.675 115.540 62.675 ;
        RECT 105.390 56.565 106.055 56.735 ;
        RECT 69.890 54.520 70.190 54.785 ;
        RECT 69.890 54.220 70.435 54.520 ;
        RECT 72.515 54.460 73.045 54.990 ;
        RECT 56.450 53.290 56.980 53.820 ;
        RECT 50.030 53.140 50.200 53.145 ;
        RECT 50.030 52.970 55.810 53.140 ;
        RECT 70.135 52.975 70.435 54.220 ;
        RECT 82.270 53.145 82.570 55.205 ;
        RECT 104.490 55.160 105.490 55.630 ;
        RECT 105.885 55.620 106.055 56.565 ;
        RECT 106.740 56.040 107.740 57.040 ;
        RECT 108.395 56.565 109.175 56.735 ;
        RECT 107.475 55.830 107.645 56.040 ;
        RECT 107.475 55.660 108.680 55.830 ;
        RECT 105.885 55.450 107.145 55.620 ;
        RECT 106.975 55.195 107.145 55.450 ;
        RECT 104.490 54.990 106.630 55.160 ;
        RECT 106.975 55.025 108.185 55.195 ;
        RECT 104.490 54.630 105.490 54.990 ;
        RECT 106.460 54.635 106.630 54.990 ;
        RECT 106.460 54.465 107.660 54.635 ;
        RECT 107.490 54.015 107.660 54.465 ;
        RECT 108.015 54.525 108.185 55.025 ;
        RECT 108.510 55.040 108.680 55.660 ;
        RECT 109.005 55.560 109.175 56.565 ;
        RECT 109.740 56.625 110.740 57.040 ;
        RECT 109.740 56.040 110.810 56.625 ;
        RECT 109.005 55.390 110.340 55.560 ;
        RECT 108.510 54.870 109.860 55.040 ;
        RECT 108.015 54.355 109.400 54.525 ;
        RECT 82.270 52.975 82.600 53.145 ;
        RECT 50.030 52.530 50.200 52.970 ;
        RECT 49.570 51.530 50.570 52.530 ;
        RECT 70.020 52.445 70.550 52.975 ;
        RECT 82.175 52.445 82.705 52.975 ;
        RECT 104.155 52.955 105.155 53.955 ;
        RECT 107.490 53.845 108.885 54.015 ;
        RECT 105.945 53.490 107.010 53.660 ;
        RECT 106.840 53.420 107.010 53.490 ;
        RECT 106.840 53.250 108.385 53.420 ;
        RECT 104.825 52.610 104.995 52.955 ;
        RECT 49.285 50.460 50.375 50.790 ;
        RECT 58.200 50.745 59.090 51.635 ;
        RECT 62.330 51.080 63.060 51.085 ;
        RECT 62.150 51.070 63.060 51.080 ;
        RECT 62.150 50.915 69.750 51.070 ;
        RECT 62.150 50.910 62.680 50.915 ;
        RECT 62.960 50.900 69.750 50.915 ;
        RECT 49.285 46.250 49.615 50.460 ;
        RECT 49.845 50.420 50.375 50.460 ;
        RECT 50.040 49.780 50.210 50.420 ;
        RECT 59.585 50.160 60.585 50.640 ;
        RECT 59.585 49.990 69.750 50.160 ;
        RECT 50.040 49.610 55.810 49.780 ;
        RECT 59.585 49.640 60.585 49.990 ;
        RECT 62.330 49.260 63.190 49.265 ;
        RECT 62.150 49.250 63.190 49.260 ;
        RECT 62.150 49.095 69.750 49.250 ;
        RECT 62.150 49.090 62.680 49.095 ;
        RECT 62.960 49.080 69.750 49.095 ;
        RECT 59.585 48.340 60.585 48.755 ;
        RECT 56.470 47.720 57.000 48.250 ;
        RECT 59.585 48.170 69.750 48.340 ;
        RECT 59.585 47.755 60.585 48.170 ;
        RECT 62.330 47.440 63.170 47.445 ;
        RECT 62.150 47.430 63.170 47.440 ;
        RECT 62.150 47.275 69.750 47.430 ;
        RECT 62.150 47.270 62.680 47.275 ;
        RECT 62.960 47.260 69.750 47.275 ;
        RECT 59.585 46.520 60.585 46.930 ;
        RECT 50.030 46.500 50.200 46.520 ;
        RECT 50.030 46.330 55.810 46.500 ;
        RECT 59.585 46.350 69.750 46.520 ;
        RECT 50.030 45.905 50.200 46.330 ;
        RECT 59.585 45.930 60.585 46.350 ;
        RECT 35.440 43.985 36.690 45.235 ;
        RECT 49.570 44.905 50.570 45.905 ;
        RECT 62.160 45.605 62.690 45.620 ;
        RECT 62.960 45.605 69.750 45.610 ;
        RECT 62.160 45.450 69.750 45.605 ;
        RECT 62.340 45.440 69.750 45.450 ;
        RECT 62.340 45.435 63.060 45.440 ;
        RECT 59.585 44.700 60.585 45.055 ;
        RECT 59.585 44.530 69.750 44.700 ;
        RECT 42.010 44.120 42.540 44.290 ;
        RECT 35.815 43.660 36.115 43.985 ;
        RECT 35.815 40.050 36.145 43.660 ;
        RECT 42.185 43.580 42.355 44.120 ;
        RECT 46.585 44.115 47.115 44.285 ;
        RECT 36.620 43.410 42.390 43.580 ;
        RECT 42.185 43.400 42.355 43.410 ;
        RECT 45.940 42.260 46.270 43.660 ;
        RECT 46.760 43.580 46.930 44.115 ;
        RECT 59.585 44.055 60.585 44.530 ;
        RECT 62.160 43.785 62.690 43.800 ;
        RECT 62.960 43.785 69.750 43.790 ;
        RECT 62.160 43.630 69.750 43.785 ;
        RECT 62.340 43.620 69.750 43.630 ;
        RECT 62.340 43.615 63.110 43.620 ;
        RECT 46.745 43.410 52.515 43.580 ;
        RECT 46.760 43.395 46.930 43.410 ;
        RECT 45.185 42.145 46.270 42.260 ;
        RECT 59.585 42.880 60.585 43.235 ;
        RECT 59.585 42.710 69.750 42.880 ;
        RECT 59.585 42.235 60.585 42.710 ;
        RECT 43.170 41.560 43.700 42.090 ;
        RECT 45.085 41.975 46.270 42.145 ;
        RECT 62.340 41.975 63.205 41.985 ;
        RECT 45.185 41.930 46.270 41.975 ;
        RECT 36.620 40.130 42.390 40.300 ;
        RECT 37.955 39.675 38.125 40.130 ;
        RECT 45.940 40.050 46.270 41.930 ;
        RECT 62.160 41.970 63.205 41.975 ;
        RECT 62.160 41.815 69.750 41.970 ;
        RECT 62.160 41.805 62.690 41.815 ;
        RECT 62.960 41.800 69.750 41.815 ;
        RECT 53.230 41.145 53.760 41.675 ;
        RECT 59.585 41.060 60.585 41.495 ;
        RECT 59.585 40.890 69.750 41.060 ;
        RECT 59.585 40.495 60.585 40.890 ;
        RECT 46.745 40.130 52.515 40.300 ;
        RECT 62.150 40.150 63.195 40.165 ;
        RECT 46.765 39.685 46.935 40.130 ;
        RECT 62.150 39.995 69.750 40.150 ;
        RECT 62.960 39.980 69.750 39.995 ;
        RECT 37.495 38.675 38.495 39.675 ;
        RECT 46.305 38.685 47.305 39.685 ;
        RECT 59.585 39.240 60.585 39.660 ;
        RECT 59.585 39.070 69.750 39.240 ;
        RECT 59.585 38.660 60.585 39.070 ;
        RECT 35.440 37.255 36.690 38.505 ;
        RECT 62.425 38.345 62.620 38.460 ;
        RECT 62.425 38.340 63.155 38.345 ;
        RECT 62.160 38.330 63.155 38.340 ;
        RECT 62.160 38.175 69.750 38.330 ;
        RECT 62.160 38.170 62.690 38.175 ;
        RECT 62.960 38.160 69.750 38.175 ;
        RECT 70.165 38.080 70.495 52.445 ;
        RECT 72.840 50.610 73.450 51.280 ;
        RECT 73.840 50.605 74.370 50.785 ;
        RECT 82.270 50.690 82.600 52.445 ;
        RECT 104.825 52.440 107.790 52.610 ;
        RECT 105.085 51.485 106.940 51.490 ;
        RECT 104.905 51.320 106.940 51.485 ;
        RECT 104.905 51.315 105.435 51.320 ;
        RECT 75.080 50.605 81.870 50.610 ;
        RECT 73.840 50.440 81.870 50.605 ;
        RECT 82.270 50.480 82.615 50.690 ;
        RECT 73.840 50.435 75.260 50.440 ;
        RECT 73.840 50.255 74.370 50.435 ;
        RECT 71.120 49.325 72.120 49.755 ;
        RECT 75.080 49.325 81.870 49.330 ;
        RECT 71.120 49.160 81.870 49.325 ;
        RECT 71.120 49.155 75.255 49.160 ;
        RECT 71.120 48.755 72.120 49.155 ;
        RECT 73.765 48.045 74.295 48.220 ;
        RECT 75.080 48.045 81.870 48.050 ;
        RECT 73.765 47.880 81.870 48.045 ;
        RECT 73.765 47.875 75.150 47.880 ;
        RECT 73.765 47.690 74.295 47.875 ;
        RECT 71.060 46.765 72.060 47.185 ;
        RECT 75.080 46.765 81.870 46.770 ;
        RECT 71.060 46.600 81.870 46.765 ;
        RECT 71.060 46.595 75.150 46.600 ;
        RECT 71.060 46.185 72.060 46.595 ;
        RECT 73.760 45.485 74.290 45.665 ;
        RECT 75.080 45.485 81.870 45.490 ;
        RECT 73.760 45.320 81.870 45.485 ;
        RECT 73.760 45.315 75.150 45.320 ;
        RECT 73.760 45.135 74.290 45.315 ;
        RECT 71.170 44.205 72.170 44.680 ;
        RECT 75.080 44.205 81.870 44.210 ;
        RECT 71.170 44.040 81.870 44.205 ;
        RECT 71.170 44.035 75.150 44.040 ;
        RECT 71.170 43.680 72.170 44.035 ;
        RECT 73.800 42.925 74.330 43.100 ;
        RECT 75.080 42.925 81.870 42.930 ;
        RECT 73.800 42.760 81.870 42.925 ;
        RECT 73.800 42.755 75.150 42.760 ;
        RECT 73.800 42.570 74.330 42.755 ;
        RECT 71.170 41.645 72.170 42.070 ;
        RECT 75.080 41.645 81.870 41.650 ;
        RECT 71.170 41.480 81.870 41.645 ;
        RECT 71.170 41.475 75.150 41.480 ;
        RECT 71.170 41.070 72.170 41.475 ;
        RECT 73.775 40.365 74.305 40.540 ;
        RECT 75.080 40.365 81.870 40.370 ;
        RECT 73.775 40.200 81.870 40.365 ;
        RECT 73.775 40.195 75.150 40.200 ;
        RECT 73.775 40.010 74.305 40.195 ;
        RECT 71.170 39.085 72.170 39.585 ;
        RECT 75.080 39.085 81.870 39.090 ;
        RECT 71.170 38.920 81.870 39.085 ;
        RECT 71.170 38.915 75.150 38.920 ;
        RECT 71.170 38.585 72.170 38.915 ;
        RECT 42.030 37.460 42.560 37.630 ;
        RECT 46.585 37.485 47.115 37.655 ;
        RECT 75.080 37.640 81.870 37.810 ;
        RECT 35.820 36.965 36.140 37.255 ;
        RECT 35.815 33.355 36.145 36.965 ;
        RECT 42.205 36.885 42.375 37.460 ;
        RECT 36.620 36.715 42.390 36.885 ;
        RECT 43.140 34.855 43.670 35.385 ;
        RECT 45.940 35.215 46.270 36.965 ;
        RECT 46.760 36.885 46.930 37.485 ;
        RECT 74.250 36.935 74.780 37.115 ;
        RECT 75.840 36.935 76.010 37.640 ;
        RECT 82.285 37.560 82.615 50.480 ;
        RECT 106.770 50.535 106.940 51.320 ;
        RECT 107.620 51.165 107.790 52.440 ;
        RECT 108.215 51.795 108.385 53.250 ;
        RECT 108.715 52.425 108.885 53.845 ;
        RECT 109.230 53.055 109.400 54.355 ;
        RECT 109.690 53.685 109.860 54.870 ;
        RECT 110.170 54.315 110.340 55.390 ;
        RECT 110.640 54.945 110.810 56.040 ;
        RECT 112.280 55.575 112.980 56.735 ;
        RECT 111.725 55.405 118.515 55.575 ;
        RECT 110.640 54.775 118.515 54.945 ;
        RECT 110.170 54.145 118.515 54.315 ;
        RECT 109.690 53.515 118.515 53.685 ;
        RECT 109.230 52.885 118.515 53.055 ;
        RECT 108.715 52.255 118.515 52.425 ;
        RECT 108.215 51.625 118.515 51.795 ;
        RECT 107.620 50.995 118.515 51.165 ;
        RECT 118.930 50.540 119.260 55.655 ;
        RECT 106.770 50.365 118.515 50.535 ;
        RECT 104.155 49.905 105.155 50.335 ;
        RECT 104.155 49.735 118.515 49.905 ;
        RECT 118.930 49.840 120.635 50.540 ;
        RECT 104.155 49.335 105.155 49.735 ;
        RECT 106.610 49.105 118.515 49.275 ;
        RECT 106.610 48.210 106.780 49.105 ;
        RECT 105.085 48.205 106.780 48.210 ;
        RECT 104.905 48.040 106.780 48.205 ;
        RECT 107.500 48.645 111.890 48.655 ;
        RECT 107.500 48.485 118.515 48.645 ;
        RECT 104.905 48.035 105.435 48.040 ;
        RECT 107.500 47.345 107.670 48.485 ;
        RECT 111.725 48.475 118.515 48.485 ;
        RECT 106.705 47.175 107.670 47.345 ;
        RECT 108.110 47.845 118.515 48.015 ;
        RECT 106.705 47.090 106.875 47.175 ;
        RECT 104.570 46.920 106.875 47.090 ;
        RECT 104.570 46.585 104.740 46.920 ;
        RECT 108.110 46.670 108.280 47.845 ;
        RECT 104.155 45.585 105.155 46.585 ;
        RECT 107.315 46.500 108.280 46.670 ;
        RECT 108.635 47.215 118.515 47.385 ;
        RECT 107.315 46.165 107.485 46.500 ;
        RECT 105.945 45.995 107.485 46.165 ;
        RECT 108.635 46.050 108.805 47.215 ;
        RECT 107.855 45.880 108.805 46.050 ;
        RECT 109.220 46.585 118.515 46.755 ;
        RECT 107.855 45.050 108.025 45.880 ;
        RECT 109.220 45.470 109.390 46.585 ;
        RECT 104.830 44.495 105.830 44.980 ;
        RECT 106.865 44.880 108.025 45.050 ;
        RECT 108.395 45.300 109.390 45.470 ;
        RECT 109.710 45.955 118.515 46.125 ;
        RECT 106.865 44.495 107.035 44.880 ;
        RECT 104.830 44.325 107.035 44.495 ;
        RECT 108.395 44.470 108.565 45.300 ;
        RECT 109.710 44.860 109.880 45.955 ;
        RECT 104.830 43.980 105.830 44.325 ;
        RECT 107.530 44.300 108.565 44.470 ;
        RECT 108.915 44.690 109.880 44.860 ;
        RECT 110.270 45.325 118.515 45.495 ;
        RECT 107.530 44.035 107.700 44.300 ;
        RECT 106.440 43.865 107.700 44.035 ;
        RECT 108.915 43.985 109.085 44.690 ;
        RECT 110.270 44.220 110.440 45.325 ;
        RECT 106.440 43.035 106.610 43.865 ;
        RECT 108.080 43.815 109.085 43.985 ;
        RECT 109.425 44.050 110.440 44.220 ;
        RECT 110.930 44.695 118.515 44.865 ;
        RECT 108.080 43.490 108.250 43.815 ;
        RECT 105.945 42.865 106.610 43.035 ;
        RECT 106.125 42.855 106.610 42.865 ;
        RECT 107.240 42.905 108.250 43.490 ;
        RECT 109.425 43.035 109.595 44.050 ;
        RECT 110.930 43.530 111.100 44.695 ;
        RECT 111.725 44.065 118.515 44.235 ;
        RECT 112.535 44.060 112.715 44.065 ;
        RECT 109.025 43.010 109.595 43.035 ;
        RECT 107.240 42.490 108.240 42.905 ;
        RECT 108.845 42.865 109.595 43.010 ;
        RECT 109.970 42.960 111.100 43.530 ;
        RECT 112.545 43.265 112.715 44.060 ;
        RECT 118.930 43.985 119.260 49.840 ;
        RECT 112.365 43.095 112.895 43.265 ;
        RECT 108.845 42.840 109.375 42.865 ;
        RECT 109.970 42.530 110.970 42.960 ;
        RECT 110.955 40.500 111.485 41.030 ;
        RECT 46.745 36.715 52.515 36.885 ;
        RECT 74.250 36.765 76.010 36.935 ;
        RECT 74.250 36.585 74.780 36.765 ;
        RECT 56.045 35.340 56.575 35.670 ;
        RECT 45.185 35.180 46.270 35.215 ;
        RECT 45.085 35.010 46.270 35.180 ;
        RECT 45.185 34.885 46.270 35.010 ;
        RECT 36.620 33.435 42.390 33.605 ;
        RECT 37.605 32.970 37.775 33.435 ;
        RECT 45.940 33.355 46.270 34.885 ;
        RECT 53.250 34.810 53.780 35.340 ;
        RECT 56.245 33.985 56.575 35.340 ;
        RECT 57.145 34.450 58.145 35.450 ;
        RECT 71.040 34.865 71.930 35.755 ;
        RECT 56.845 33.985 57.175 34.030 ;
        RECT 56.245 33.655 57.175 33.985 ;
        RECT 57.645 33.950 57.815 34.450 ;
        RECT 57.590 33.780 64.380 33.950 ;
        RECT 46.745 33.435 52.515 33.605 ;
        RECT 46.750 32.980 46.920 33.435 ;
        RECT 35.440 31.160 36.690 32.410 ;
        RECT 37.145 31.970 38.145 32.970 ;
        RECT 46.290 31.980 47.290 32.980 ;
        RECT 56.845 32.790 57.175 33.655 ;
        RECT 64.750 33.090 65.360 33.760 ;
        RECT 70.295 33.735 70.625 34.205 ;
        RECT 71.475 34.125 71.645 34.865 ;
        RECT 71.040 33.955 77.830 34.125 ;
        RECT 69.225 33.675 70.625 33.735 ;
        RECT 69.125 33.505 70.625 33.675 ;
        RECT 69.225 33.405 70.625 33.505 ;
        RECT 57.590 32.870 64.380 33.040 ;
        RECT 70.295 32.965 70.625 33.405 ;
        RECT 71.040 33.045 77.830 33.215 ;
        RECT 78.800 33.210 79.410 33.880 ;
        RECT 57.605 32.405 57.775 32.870 ;
        RECT 41.990 31.345 42.520 31.515 ;
        RECT 35.825 30.850 36.145 31.160 ;
        RECT 35.815 27.240 36.145 30.850 ;
        RECT 42.165 30.770 42.335 31.345 ;
        RECT 47.775 31.325 48.305 31.495 ;
        RECT 57.145 31.405 58.145 32.405 ;
        RECT 71.685 32.325 71.855 33.045 ;
        RECT 71.505 31.795 72.035 32.325 ;
        RECT 36.620 30.600 42.390 30.770 ;
        RECT 43.140 28.765 43.670 29.295 ;
        RECT 45.940 28.975 46.270 30.850 ;
        RECT 47.950 30.770 48.120 31.325 ;
        RECT 46.745 30.600 52.515 30.770 ;
        RECT 45.085 28.645 46.270 28.975 ;
        RECT 53.250 28.785 53.780 29.315 ;
        RECT 36.620 27.320 42.390 27.490 ;
        RECT 37.605 26.855 37.775 27.320 ;
        RECT 45.940 27.240 46.270 28.645 ;
        RECT 46.785 27.490 46.955 27.500 ;
        RECT 46.745 27.320 52.515 27.490 ;
        RECT 46.785 26.885 46.955 27.320 ;
        RECT 35.610 24.790 36.860 26.040 ;
        RECT 37.145 25.855 38.145 26.855 ;
        RECT 46.325 25.885 47.325 26.885 ;
        RECT 61.705 26.405 61.875 27.075 ;
        RECT 42.030 24.920 42.560 25.090 ;
        RECT 47.775 24.920 48.305 25.090 ;
        RECT 35.830 24.445 36.130 24.790 ;
        RECT 35.815 20.835 36.145 24.445 ;
        RECT 42.205 24.365 42.375 24.920 ;
        RECT 36.620 24.195 42.390 24.365 ;
        RECT 45.940 22.890 46.270 24.445 ;
        RECT 47.950 24.365 48.120 24.920 ;
        RECT 46.745 24.195 52.515 24.365 ;
        RECT 61.705 23.985 61.875 25.865 ;
        RECT 86.770 25.195 86.940 27.075 ;
        RECT 45.185 22.820 46.270 22.890 ;
        RECT 43.140 22.290 43.670 22.820 ;
        RECT 45.085 22.650 46.270 22.820 ;
        RECT 45.185 22.560 46.270 22.650 ;
        RECT 36.620 21.075 42.390 21.085 ;
        RECT 36.615 20.915 42.390 21.075 ;
        RECT 36.615 20.460 36.785 20.915 ;
        RECT 45.940 20.835 46.270 22.560 ;
        RECT 53.250 22.440 53.780 22.970 ;
        RECT 61.705 21.565 61.875 23.445 ;
        RECT 86.770 22.775 86.940 24.655 ;
        RECT 86.770 21.565 86.940 22.235 ;
        RECT 46.740 21.085 46.910 21.095 ;
        RECT 46.740 20.915 52.515 21.085 ;
        RECT 46.740 20.480 46.910 20.915 ;
        RECT 36.155 19.460 37.155 20.460 ;
        RECT 46.280 19.480 47.280 20.480 ;
      LAYER met1 ;
        RECT 85.970 220.725 86.970 220.820 ;
        RECT 9.315 219.725 86.970 220.725 ;
        RECT 9.315 3.005 10.315 219.725 ;
        RECT 61.085 218.925 62.085 219.725 ;
        RECT 85.970 218.925 86.970 219.725 ;
        RECT 37.665 213.285 43.340 218.925 ;
        RECT 56.285 213.425 66.285 218.925 ;
        RECT 84.025 213.515 94.025 218.925 ;
        RECT 95.740 216.635 114.670 217.335 ;
        RECT 37.665 212.585 54.495 213.285 ;
        RECT 37.665 188.830 43.340 212.585 ;
        RECT 51.710 211.265 52.410 212.585 ;
        RECT 51.710 210.565 52.465 211.265 ;
        RECT 51.730 208.220 52.430 210.565 ;
        RECT 58.980 210.360 59.570 211.010 ;
        RECT 53.505 208.640 54.095 209.290 ;
        RECT 51.730 207.520 54.485 208.220 ;
        RECT 51.730 206.365 52.430 207.520 ;
        RECT 51.730 205.665 52.465 206.365 ;
        RECT 59.125 206.355 59.425 210.360 ;
        RECT 62.665 208.870 63.365 213.425 ;
        RECT 64.080 209.570 64.670 210.220 ;
        RECT 91.575 208.870 92.275 213.515 ;
        RECT 93.165 209.570 93.755 210.220 ;
        RECT 62.540 207.860 63.490 208.870 ;
        RECT 91.450 207.860 92.400 208.870 ;
        RECT 58.980 205.705 59.570 206.355 ;
        RECT 63.900 205.765 64.490 206.415 ;
        RECT 93.165 205.785 93.755 206.435 ;
        RECT 51.750 201.790 52.450 205.665 ;
        RECT 53.465 203.830 54.055 204.480 ;
        RECT 51.750 201.090 54.410 201.790 ;
        RECT 51.750 199.130 52.505 201.090 ;
        RECT 59.125 199.960 59.425 205.705 ;
        RECT 95.740 205.475 96.440 216.635 ;
        RECT 98.965 216.045 99.555 216.220 ;
        RECT 93.920 205.460 96.440 205.475 ;
        RECT 63.905 204.655 64.485 205.295 ;
        RECT 65.120 204.775 96.440 205.460 ;
        RECT 96.880 215.745 99.555 216.045 ;
        RECT 96.880 208.850 97.180 215.745 ;
        RECT 98.965 215.570 99.555 215.745 ;
        RECT 104.590 214.765 105.190 216.635 ;
        RECT 107.245 215.965 107.835 216.220 ;
        RECT 104.575 214.115 105.190 214.765 ;
        RECT 97.600 212.950 98.200 213.590 ;
        RECT 103.030 209.780 103.620 210.430 ;
        RECT 98.965 208.850 99.555 209.025 ;
        RECT 96.880 208.550 99.555 208.850 ;
        RECT 65.120 204.760 94.620 204.775 ;
        RECT 65.120 204.690 65.820 204.760 ;
        RECT 58.980 199.310 59.570 199.960 ;
        RECT 51.750 196.865 52.450 199.130 ;
        RECT 53.520 197.885 54.110 198.060 ;
        RECT 59.125 197.885 59.425 199.310 ;
        RECT 53.520 197.585 59.425 197.885 ;
        RECT 53.520 197.410 54.110 197.585 ;
        RECT 51.750 196.165 54.465 196.865 ;
        RECT 51.750 195.140 52.450 196.165 ;
        RECT 51.750 194.440 52.465 195.140 ;
        RECT 59.125 194.915 59.425 197.585 ;
        RECT 58.980 194.265 59.570 194.915 ;
        RECT 53.520 193.065 54.110 193.240 ;
        RECT 59.125 193.065 59.425 194.265 ;
        RECT 53.520 192.765 59.425 193.065 ;
        RECT 53.520 192.590 54.110 192.765 ;
        RECT 53.665 190.310 53.965 192.590 ;
        RECT 53.455 189.670 54.035 190.310 ;
        RECT 37.665 188.780 47.285 188.830 ;
        RECT 37.665 188.130 55.865 188.780 ;
        RECT 37.665 184.100 43.340 188.130 ;
        RECT 44.570 186.870 45.270 188.130 ;
        RECT 46.585 188.080 55.865 188.130 ;
        RECT 53.840 185.995 54.430 186.645 ;
        RECT 52.830 184.645 53.420 184.820 ;
        RECT 53.985 184.645 54.285 185.995 ;
        RECT 54.445 184.645 55.025 184.810 ;
        RECT 52.830 184.345 55.025 184.645 ;
        RECT 52.830 184.170 53.420 184.345 ;
        RECT 37.665 183.400 47.230 184.100 ;
        RECT 37.665 179.525 43.340 183.400 ;
        RECT 44.560 182.415 45.260 183.400 ;
        RECT 53.985 182.190 54.285 184.345 ;
        RECT 54.445 184.170 55.025 184.345 ;
        RECT 53.840 181.540 54.430 182.190 ;
        RECT 52.830 180.130 53.420 180.305 ;
        RECT 53.985 180.130 54.285 181.540 ;
        RECT 52.830 179.830 54.285 180.130 ;
        RECT 52.830 179.655 53.420 179.830 ;
        RECT 37.665 179.510 47.120 179.525 ;
        RECT 37.665 178.860 47.230 179.510 ;
        RECT 37.665 178.825 47.120 178.860 ;
        RECT 37.665 173.985 43.340 178.825 ;
        RECT 44.560 177.815 45.260 178.825 ;
        RECT 53.985 177.495 54.285 179.830 ;
        RECT 55.165 178.415 55.865 188.080 ;
        RECT 56.630 186.985 57.210 187.160 ;
        RECT 64.045 186.985 64.345 204.655 ;
        RECT 83.300 203.160 84.000 204.760 ;
        RECT 81.530 202.460 84.000 203.160 ;
        RECT 76.220 200.365 76.800 201.005 ;
        RECT 76.380 199.975 76.680 200.365 ;
        RECT 76.245 199.325 76.835 199.975 ;
        RECT 76.380 196.905 76.680 199.325 ;
        RECT 77.690 196.905 78.280 197.080 ;
        RECT 76.380 196.605 78.280 196.905 ;
        RECT 76.380 192.700 76.680 196.605 ;
        RECT 77.690 196.430 78.280 196.605 ;
        RECT 83.300 196.055 84.000 202.460 ;
        RECT 81.530 195.355 84.000 196.055 ;
        RECT 83.300 194.255 84.000 195.355 ;
        RECT 96.880 201.875 97.180 208.550 ;
        RECT 98.965 208.375 99.555 208.550 ;
        RECT 97.600 205.775 98.200 206.415 ;
        RECT 103.115 202.715 103.705 203.365 ;
        RECT 98.965 201.875 99.555 202.050 ;
        RECT 96.880 201.575 99.555 201.875 ;
        RECT 96.880 194.865 97.180 201.575 ;
        RECT 98.965 201.400 99.555 201.575 ;
        RECT 97.600 198.825 98.200 199.465 ;
        RECT 103.115 195.835 103.705 196.485 ;
        RECT 98.965 194.865 99.555 195.075 ;
        RECT 96.880 194.565 99.555 194.865 ;
        RECT 76.225 192.050 76.815 192.700 ;
        RECT 76.370 190.075 76.670 192.050 ;
        RECT 95.830 191.750 96.430 192.390 ;
        RECT 77.690 190.075 78.280 190.215 ;
        RECT 76.370 189.775 78.280 190.075 ;
        RECT 76.370 188.960 76.670 189.775 ;
        RECT 77.690 189.565 78.280 189.775 ;
        RECT 95.980 188.960 96.280 191.750 ;
        RECT 76.370 188.660 96.280 188.960 ;
        RECT 76.370 188.655 76.670 188.660 ;
        RECT 96.880 187.980 97.180 194.565 ;
        RECT 98.965 194.425 99.555 194.565 ;
        RECT 104.590 192.585 105.190 214.115 ;
        RECT 105.460 215.825 107.835 215.965 ;
        RECT 105.460 208.770 105.600 215.825 ;
        RECT 107.245 215.570 107.835 215.825 ;
        RECT 113.970 214.640 114.670 216.635 ;
        RECT 112.675 213.940 114.670 214.640 ;
        RECT 105.795 213.090 106.395 213.730 ;
        RECT 106.950 209.780 107.540 210.430 ;
        RECT 107.245 208.770 107.835 209.025 ;
        RECT 105.460 208.630 107.835 208.770 ;
        RECT 105.460 201.865 105.600 208.630 ;
        RECT 107.245 208.375 107.835 208.630 ;
        RECT 113.970 207.875 114.670 213.940 ;
        RECT 112.675 207.175 114.670 207.875 ;
        RECT 105.795 206.010 106.395 206.650 ;
        RECT 107.035 202.715 107.625 203.365 ;
        RECT 107.245 201.865 107.835 202.120 ;
        RECT 105.460 201.725 107.835 201.865 ;
        RECT 105.460 194.885 105.600 201.725 ;
        RECT 107.245 201.470 107.835 201.725 ;
        RECT 112.620 200.680 113.320 200.740 ;
        RECT 113.970 200.680 114.670 207.175 ;
        RECT 112.620 199.980 114.670 200.680 ;
        RECT 105.795 199.140 106.395 199.780 ;
        RECT 107.035 195.835 107.625 196.485 ;
        RECT 107.245 194.885 107.835 195.140 ;
        RECT 105.460 194.745 107.835 194.885 ;
        RECT 97.600 191.800 98.200 192.440 ;
        RECT 103.115 188.675 103.705 189.325 ;
        RECT 105.460 187.980 105.600 194.745 ;
        RECT 107.245 194.490 107.835 194.745 ;
        RECT 113.970 193.260 114.670 199.980 ;
        RECT 120.160 193.260 124.665 218.925 ;
        RECT 112.675 192.560 124.665 193.260 ;
        RECT 105.795 191.800 106.395 192.440 ;
        RECT 107.035 188.675 107.625 189.325 ;
        RECT 96.880 187.680 119.740 187.980 ;
        RECT 56.630 186.685 64.345 186.985 ;
        RECT 56.630 186.520 57.210 186.685 ;
        RECT 58.525 184.050 58.755 185.910 ;
        RECT 118.860 185.710 119.090 185.910 ;
        RECT 119.440 185.710 119.740 187.680 ;
        RECT 118.860 185.570 119.740 185.710 ;
        RECT 118.860 185.260 119.090 185.570 ;
        RECT 58.525 181.630 58.755 183.490 ;
        RECT 118.860 182.840 119.090 184.700 ;
        RECT 58.525 179.210 58.755 181.070 ;
        RECT 118.860 180.420 119.090 182.280 ;
        RECT 120.160 179.860 124.665 192.560 ;
        RECT 118.860 179.210 124.665 179.860 ;
        RECT 55.165 177.715 88.700 178.415 ;
        RECT 53.840 176.845 54.430 177.495 ;
        RECT 52.830 175.525 53.420 175.705 ;
        RECT 53.985 175.525 54.285 176.845 ;
        RECT 52.830 175.225 54.285 175.525 ;
        RECT 52.830 175.055 53.420 175.225 ;
        RECT 37.665 173.940 46.720 173.985 ;
        RECT 37.665 173.290 47.145 173.940 ;
        RECT 37.665 173.285 46.720 173.290 ;
        RECT 37.665 169.505 43.340 173.285 ;
        RECT 44.560 172.270 45.260 173.285 ;
        RECT 53.985 171.785 54.285 175.225 ;
        RECT 88.000 174.560 88.700 177.715 ;
        RECT 104.890 176.215 113.745 176.915 ;
        RECT 89.230 175.555 89.820 176.205 ;
        RECT 87.875 173.550 88.825 174.560 ;
        RECT 104.890 174.290 105.590 176.215 ;
        RECT 107.065 176.045 107.655 176.215 ;
        RECT 91.170 173.590 105.590 174.290 ;
        RECT 113.045 174.955 113.745 176.215 ;
        RECT 120.160 174.955 124.665 179.210 ;
        RECT 113.045 174.255 124.665 174.955 ;
        RECT 53.815 171.135 54.405 171.785 ;
        RECT 37.665 168.805 47.200 169.505 ;
        RECT 52.595 169.455 53.185 170.105 ;
        RECT 37.665 164.850 43.340 168.805 ;
        RECT 44.640 167.655 45.340 168.805 ;
        RECT 53.985 167.475 54.285 171.135 ;
        RECT 53.845 166.825 54.435 167.475 ;
        RECT 46.500 164.850 47.200 164.915 ;
        RECT 37.665 164.150 47.200 164.850 ;
        RECT 52.530 164.820 53.120 165.470 ;
        RECT 21.395 148.670 23.635 148.735 ;
        RECT 37.665 148.670 43.340 164.150 ;
        RECT 44.560 163.165 45.260 164.150 ;
        RECT 53.985 162.875 54.285 166.825 ;
        RECT 88.000 164.600 88.700 173.550 ;
        RECT 89.255 171.585 89.845 172.235 ;
        RECT 89.245 165.495 89.835 166.145 ;
        RECT 87.965 163.590 88.915 164.600 ;
        RECT 92.280 164.370 92.980 173.590 ;
        RECT 105.765 172.735 106.365 173.375 ;
        RECT 107.285 170.780 107.875 170.870 ;
        RECT 105.165 170.480 107.875 170.780 ;
        RECT 93.970 165.960 94.560 166.175 ;
        RECT 105.165 165.960 105.465 170.480 ;
        RECT 107.285 170.220 107.875 170.480 ;
        RECT 107.010 169.470 107.710 169.525 ;
        RECT 107.010 168.770 113.735 169.470 ;
        RECT 113.035 168.400 113.735 168.770 ;
        RECT 120.160 168.400 124.665 174.255 ;
        RECT 113.035 167.725 124.665 168.400 ;
        RECT 113.090 167.700 124.665 167.725 ;
        RECT 93.970 165.660 105.465 165.960 ;
        RECT 105.765 165.945 106.365 166.585 ;
        RECT 93.970 165.525 94.560 165.660 ;
        RECT 91.180 163.670 92.980 164.370 ;
        RECT 105.165 163.565 105.465 165.660 ;
        RECT 107.285 163.565 107.875 163.740 ;
        RECT 105.165 163.265 107.875 163.565 ;
        RECT 107.285 163.090 107.875 163.265 ;
        RECT 53.825 162.225 54.415 162.875 ;
        RECT 86.115 162.085 86.730 162.090 ;
        RECT 86.080 160.720 86.730 162.085 ;
        RECT 89.255 161.595 89.845 162.245 ;
        RECT 52.535 160.070 53.125 160.720 ;
        RECT 55.475 160.020 113.620 160.720 ;
        RECT 86.080 160.010 86.730 160.020 ;
        RECT 112.920 158.250 113.620 160.020 ;
        RECT 45.885 156.390 46.115 158.250 ;
        RECT 110.890 157.600 113.620 158.250 ;
        RECT 45.885 153.970 46.115 155.830 ;
        RECT 110.890 155.180 111.120 157.040 ;
        RECT 45.885 151.550 46.115 153.410 ;
        RECT 110.890 152.760 111.120 154.620 ;
        RECT 45.885 149.130 46.115 150.990 ;
        RECT 110.890 150.340 111.120 152.200 ;
        RECT 21.395 146.670 43.340 148.670 ;
        RECT 45.885 146.710 46.115 148.570 ;
        RECT 110.890 147.920 111.120 149.780 ;
        RECT 21.395 146.535 23.635 146.670 ;
        RECT 37.665 138.890 43.340 146.670 ;
        RECT 45.885 144.290 46.115 146.150 ;
        RECT 110.890 145.500 111.120 147.360 ;
        RECT 112.920 145.825 113.620 157.600 ;
        RECT 120.160 147.670 124.665 167.700 ;
        RECT 138.245 147.670 140.485 147.750 ;
        RECT 45.885 141.870 46.115 143.730 ;
        RECT 110.890 143.080 111.120 144.940 ;
        RECT 45.885 139.450 46.115 141.310 ;
        RECT 110.890 140.660 111.120 142.520 ;
        RECT 110.890 139.450 112.190 140.100 ;
        RECT 111.540 138.890 112.190 139.450 ;
        RECT 37.665 138.240 112.190 138.890 ;
        RECT 37.665 137.925 43.340 138.240 ;
        RECT 112.665 137.925 117.665 145.825 ;
        RECT 120.160 145.670 140.485 147.670 ;
        RECT 120.160 137.925 124.665 145.670 ;
        RECT 138.245 145.550 140.485 145.670 ;
        RECT 114.655 115.400 115.655 137.925 ;
        RECT 14.125 114.400 115.655 115.400 ;
        RECT 14.125 4.480 15.125 114.400 ;
        RECT 28.785 88.175 34.895 110.390 ;
        RECT 44.050 108.140 44.950 108.300 ;
        RECT 53.035 108.150 53.935 108.310 ;
        RECT 63.270 108.150 64.170 108.310 ;
        RECT 44.030 107.500 44.970 108.140 ;
        RECT 53.015 107.510 53.955 108.150 ;
        RECT 63.250 107.510 64.190 108.150 ;
        RECT 71.675 108.125 72.255 108.765 ;
        RECT 76.775 108.675 77.675 108.835 ;
        RECT 44.050 107.340 44.950 107.500 ;
        RECT 53.035 107.350 53.935 107.510 ;
        RECT 63.270 107.350 64.170 107.510 ;
        RECT 42.295 105.625 43.195 105.785 ;
        RECT 42.275 104.985 43.215 105.625 ;
        RECT 59.510 105.480 60.410 105.640 ;
        RECT 69.535 105.480 70.435 105.640 ;
        RECT 42.295 104.825 43.195 104.985 ;
        RECT 49.745 104.690 50.335 105.340 ;
        RECT 59.490 104.840 60.430 105.480 ;
        RECT 69.515 104.840 70.455 105.480 ;
        RECT 71.785 105.135 71.925 108.125 ;
        RECT 76.755 108.035 77.695 108.675 ;
        RECT 76.775 107.875 77.675 108.035 ;
        RECT 79.960 106.560 80.540 106.745 ;
        RECT 124.160 106.560 129.040 110.390 ;
        RECT 79.915 105.860 129.040 106.560 ;
        RECT 43.975 101.155 44.975 102.155 ;
        RECT 44.050 99.290 44.950 99.450 ;
        RECT 44.030 98.650 44.970 99.290 ;
        RECT 44.050 98.490 44.950 98.650 ;
        RECT 49.985 96.465 50.125 104.690 ;
        RECT 59.510 104.680 60.410 104.840 ;
        RECT 69.535 104.680 70.435 104.840 ;
        RECT 71.545 104.485 72.135 105.135 ;
        RECT 80.365 104.855 80.945 105.050 ;
        RECT 80.365 104.715 81.315 104.855 ;
        RECT 52.185 102.725 52.775 103.375 ;
        RECT 49.970 96.265 50.125 96.465 ;
        RECT 42.295 95.830 43.195 95.990 ;
        RECT 42.275 95.190 43.215 95.830 ;
        RECT 49.970 95.230 50.110 96.265 ;
        RECT 42.295 95.030 43.195 95.190 ;
        RECT 49.765 94.580 50.355 95.230 ;
        RECT 43.975 91.245 44.975 92.245 ;
        RECT 35.375 88.175 35.955 88.425 ;
        RECT 28.785 88.035 35.955 88.175 ;
        RECT 44.050 88.070 44.950 88.230 ;
        RECT 28.785 57.180 34.895 88.035 ;
        RECT 35.375 87.785 35.955 88.035 ;
        RECT 44.030 87.430 44.970 88.070 ;
        RECT 44.050 87.270 44.950 87.430 ;
        RECT 42.295 86.470 43.195 86.630 ;
        RECT 42.275 85.830 43.215 86.470 ;
        RECT 42.295 85.670 43.195 85.830 ;
        RECT 49.970 85.155 50.110 94.580 ;
        RECT 52.410 93.445 52.550 102.725 ;
        RECT 62.345 102.695 62.935 103.345 ;
        RECT 52.960 101.190 53.960 102.190 ;
        RECT 62.565 99.015 62.705 102.695 ;
        RECT 63.455 101.130 64.455 102.130 ;
        RECT 71.785 101.800 71.925 104.485 ;
        RECT 80.365 104.410 80.945 104.715 ;
        RECT 81.175 103.910 81.315 104.715 ;
        RECT 81.120 103.260 81.350 103.910 ;
        RECT 72.395 101.800 73.345 102.170 ;
        RECT 71.785 101.660 73.345 101.800 ;
        RECT 77.425 101.765 78.325 101.925 ;
        RECT 71.785 99.015 71.925 101.660 ;
        RECT 72.395 101.160 73.345 101.660 ;
        RECT 77.405 101.125 78.345 101.765 ;
        RECT 77.425 100.965 78.325 101.125 ;
        RECT 81.120 100.840 81.350 102.700 ;
        RECT 121.955 102.050 122.185 103.910 ;
        RECT 62.565 98.875 71.925 99.015 ;
        RECT 53.035 98.190 53.935 98.350 ;
        RECT 53.015 97.550 53.955 98.190 ;
        RECT 53.035 97.390 53.935 97.550 ;
        RECT 62.565 97.150 62.705 98.875 ;
        RECT 63.270 98.210 64.170 98.370 ;
        RECT 63.250 97.570 64.190 98.210 ;
        RECT 63.270 97.410 64.170 97.570 ;
        RECT 62.345 96.500 62.935 97.150 ;
        RECT 59.510 95.130 60.410 95.290 ;
        RECT 59.490 94.490 60.430 95.130 ;
        RECT 59.510 94.330 60.410 94.490 ;
        RECT 52.185 92.795 52.775 93.445 ;
        RECT 49.745 84.505 50.335 85.155 ;
        RECT 43.975 81.090 44.975 82.090 ;
        RECT 44.050 78.995 44.950 79.155 ;
        RECT 44.030 78.355 44.970 78.995 ;
        RECT 44.050 78.195 44.950 78.355 ;
        RECT 41.690 75.985 42.590 76.145 ;
        RECT 41.670 75.345 42.610 75.985 ;
        RECT 49.970 75.955 50.110 84.505 ;
        RECT 52.410 83.395 52.550 92.795 ;
        RECT 52.960 91.280 53.960 92.280 ;
        RECT 53.035 88.420 53.935 88.580 ;
        RECT 53.015 87.780 53.955 88.420 ;
        RECT 53.035 87.620 53.935 87.780 ;
        RECT 62.565 87.145 62.705 96.500 ;
        RECT 69.535 95.130 70.435 95.290 ;
        RECT 71.785 95.170 71.925 98.875 ;
        RECT 76.700 98.675 77.600 98.835 ;
        RECT 76.680 98.035 77.620 98.675 ;
        RECT 81.120 98.420 81.350 100.280 ;
        RECT 121.955 99.630 122.185 101.490 ;
        RECT 124.160 99.075 129.040 105.860 ;
        RECT 122.080 99.070 129.040 99.075 ;
        RECT 121.955 98.420 129.040 99.070 ;
        RECT 122.080 98.375 129.040 98.420 ;
        RECT 76.700 97.875 77.600 98.035 ;
        RECT 124.160 97.875 129.040 98.375 ;
        RECT 120.200 97.175 129.040 97.875 ;
        RECT 91.525 96.700 110.835 96.840 ;
        RECT 69.515 94.490 70.455 95.130 ;
        RECT 71.565 94.520 72.155 95.170 ;
        RECT 91.525 95.110 91.665 96.700 ;
        RECT 110.695 95.705 110.835 96.700 ;
        RECT 91.410 94.840 92.000 95.110 ;
        RECT 84.245 94.700 92.000 94.840 ;
        RECT 69.535 94.330 70.435 94.490 ;
        RECT 63.455 91.235 64.455 92.235 ;
        RECT 71.785 91.790 71.925 94.520 ;
        RECT 72.395 91.790 73.345 92.270 ;
        RECT 77.425 92.245 78.325 92.405 ;
        RECT 71.785 91.650 73.345 91.790 ;
        RECT 63.270 88.545 64.170 88.705 ;
        RECT 63.250 87.905 64.190 88.545 ;
        RECT 63.270 87.745 64.170 87.905 ;
        RECT 62.345 86.495 62.935 87.145 ;
        RECT 59.510 85.110 60.410 85.270 ;
        RECT 59.490 84.470 60.430 85.110 ;
        RECT 59.510 84.310 60.410 84.470 ;
        RECT 52.185 82.745 52.775 83.395 ;
        RECT 52.400 79.805 52.540 82.745 ;
        RECT 52.960 81.265 53.960 82.265 ;
        RECT 62.570 79.805 62.710 86.495 ;
        RECT 69.535 85.270 70.435 85.430 ;
        RECT 71.785 85.410 71.925 91.650 ;
        RECT 72.395 91.260 73.345 91.650 ;
        RECT 77.405 91.605 78.345 92.245 ;
        RECT 77.425 91.445 78.325 91.605 ;
        RECT 76.700 88.845 77.600 89.005 ;
        RECT 76.680 88.205 77.620 88.845 ;
        RECT 76.700 88.045 77.600 88.205 ;
        RECT 69.515 84.630 70.455 85.270 ;
        RECT 71.505 84.760 72.095 85.410 ;
        RECT 69.535 84.470 70.435 84.630 ;
        RECT 71.785 83.505 71.925 84.760 ;
        RECT 71.770 83.365 71.925 83.505 ;
        RECT 63.455 81.380 64.455 82.380 ;
        RECT 52.400 79.665 62.710 79.805 ;
        RECT 52.400 77.975 52.540 79.665 ;
        RECT 53.035 78.985 53.935 79.145 ;
        RECT 53.015 78.345 53.955 78.985 ;
        RECT 53.035 78.185 53.935 78.345 ;
        RECT 52.185 77.325 52.775 77.975 ;
        RECT 62.570 77.880 62.710 79.665 ;
        RECT 63.270 79.030 64.170 79.190 ;
        RECT 63.250 78.390 64.190 79.030 ;
        RECT 63.270 78.230 64.170 78.390 ;
        RECT 62.345 77.230 62.935 77.880 ;
        RECT 59.510 76.175 60.410 76.335 ;
        RECT 49.765 75.690 50.355 75.955 ;
        RECT 50.540 75.690 51.120 75.940 ;
        RECT 49.765 75.550 51.120 75.690 ;
        RECT 41.690 75.185 42.590 75.345 ;
        RECT 49.765 75.305 50.355 75.550 ;
        RECT 50.540 75.300 51.120 75.550 ;
        RECT 59.490 75.535 60.430 76.175 ;
        RECT 69.535 75.945 70.435 76.105 ;
        RECT 59.510 75.375 60.410 75.535 ;
        RECT 69.515 75.305 70.455 75.945 ;
        RECT 71.785 75.710 71.925 83.365 ;
        RECT 72.500 81.530 73.500 82.530 ;
        RECT 77.390 81.890 78.290 82.050 ;
        RECT 77.370 81.250 78.310 81.890 ;
        RECT 77.390 81.090 78.290 81.250 ;
        RECT 76.860 78.720 77.760 78.880 ;
        RECT 76.840 78.080 77.780 78.720 ;
        RECT 76.860 77.920 77.760 78.080 ;
        RECT 84.245 76.095 84.385 94.700 ;
        RECT 91.410 94.460 92.000 94.700 ;
        RECT 94.645 94.455 95.645 95.455 ;
        RECT 96.150 95.080 97.050 95.240 ;
        RECT 96.130 94.440 97.070 95.080 ;
        RECT 110.445 95.055 111.035 95.705 ;
        RECT 112.975 94.455 113.975 95.455 ;
        RECT 114.480 95.080 115.380 95.240 ;
        RECT 114.460 94.440 115.400 95.080 ;
        RECT 96.150 94.280 97.050 94.440 ;
        RECT 114.480 94.280 115.380 94.440 ;
        RECT 94.220 93.830 95.120 93.990 ;
        RECT 112.550 93.830 113.450 93.990 ;
        RECT 92.740 92.730 93.740 93.730 ;
        RECT 94.200 93.190 95.140 93.830 ;
        RECT 94.220 93.030 95.120 93.190 ;
        RECT 91.710 91.165 92.710 92.165 ;
        RECT 93.170 92.160 94.070 92.320 ;
        RECT 93.150 91.520 94.090 92.160 ;
        RECT 102.775 92.045 103.775 93.045 ;
        RECT 111.070 92.730 112.070 93.730 ;
        RECT 112.530 93.190 113.470 93.830 ;
        RECT 112.550 93.030 113.450 93.190 ;
        RECT 93.170 91.360 94.070 91.520 ;
        RECT 110.040 91.165 111.040 92.165 ;
        RECT 111.500 92.160 112.400 92.320 ;
        RECT 111.480 91.520 112.420 92.160 ;
        RECT 111.500 91.360 112.400 91.520 ;
        RECT 87.855 89.765 88.755 89.925 ;
        RECT 87.835 89.125 88.775 89.765 ;
        RECT 89.360 89.660 90.360 90.660 ;
        RECT 91.055 90.580 91.955 90.740 ;
        RECT 91.035 89.940 91.975 90.580 ;
        RECT 91.055 89.780 91.955 89.940 ;
        RECT 106.185 89.765 107.085 89.925 ;
        RECT 106.165 89.125 107.105 89.765 ;
        RECT 107.690 89.660 108.690 90.660 ;
        RECT 109.385 90.580 110.285 90.740 ;
        RECT 109.365 89.940 110.305 90.580 ;
        RECT 109.385 89.780 110.285 89.940 ;
        RECT 87.855 88.965 88.755 89.125 ;
        RECT 106.185 88.965 107.085 89.125 ;
        RECT 86.145 87.500 87.145 88.500 ;
        RECT 87.855 87.405 88.755 87.565 ;
        RECT 104.475 87.520 105.475 88.520 ;
        RECT 124.160 88.475 129.040 97.175 ;
        RECT 120.065 87.775 129.040 88.475 ;
        RECT 106.185 87.405 107.085 87.565 ;
        RECT 87.835 86.765 88.775 87.405 ;
        RECT 106.165 86.765 107.105 87.405 ;
        RECT 87.855 86.605 88.755 86.765 ;
        RECT 106.185 86.605 107.085 86.765 ;
        RECT 88.680 85.120 89.680 86.120 ;
        RECT 90.190 85.940 91.090 86.100 ;
        RECT 90.170 85.300 91.110 85.940 ;
        RECT 90.190 85.140 91.090 85.300 ;
        RECT 107.010 85.120 108.010 86.120 ;
        RECT 108.520 85.940 109.420 86.100 ;
        RECT 108.500 85.300 109.440 85.940 ;
        RECT 108.520 85.140 109.420 85.300 ;
        RECT 90.755 83.695 91.755 84.695 ;
        RECT 92.295 84.420 93.195 84.580 ;
        RECT 92.275 83.780 93.215 84.420 ;
        RECT 92.295 83.620 93.195 83.780 ;
        RECT 109.085 83.695 110.085 84.695 ;
        RECT 110.625 84.420 111.525 84.580 ;
        RECT 110.605 83.780 111.545 84.420 ;
        RECT 110.625 83.620 111.525 83.780 ;
        RECT 90.755 81.750 91.755 82.750 ;
        RECT 92.500 82.595 93.400 82.755 ;
        RECT 92.480 81.955 93.420 82.595 ;
        RECT 92.500 81.795 93.400 81.955 ;
        RECT 109.085 81.750 110.085 82.750 ;
        RECT 110.830 82.595 111.730 82.755 ;
        RECT 110.810 81.955 111.750 82.595 ;
        RECT 110.830 81.795 111.730 81.955 ;
        RECT 93.025 80.210 94.025 81.210 ;
        RECT 94.580 81.135 95.480 81.295 ;
        RECT 94.560 80.495 95.500 81.135 ;
        RECT 94.580 80.335 95.480 80.495 ;
        RECT 96.180 80.210 97.180 81.210 ;
        RECT 111.355 80.210 112.355 81.210 ;
        RECT 112.910 81.135 113.810 81.295 ;
        RECT 112.890 80.495 113.830 81.135 ;
        RECT 112.910 80.335 113.810 80.495 ;
        RECT 114.510 80.210 115.510 81.210 ;
        RECT 91.275 77.860 110.115 78.000 ;
        RECT 91.275 76.725 91.415 77.860 ;
        RECT 91.100 76.095 91.690 76.725 ;
        RECT 94.405 76.165 95.405 77.165 ;
        RECT 95.860 76.790 96.760 76.950 ;
        RECT 95.840 76.150 96.780 76.790 ;
        RECT 109.975 76.350 110.115 77.860 ;
        RECT 84.245 76.075 91.690 76.095 ;
        RECT 84.245 75.955 91.415 76.075 ;
        RECT 95.860 75.990 96.760 76.150 ;
        RECT 69.535 75.145 70.435 75.305 ;
        RECT 71.525 75.060 72.115 75.710 ;
        RECT 43.975 72.085 44.975 73.085 ;
        RECT 52.960 72.060 53.960 73.060 ;
        RECT 63.455 72.205 64.455 73.205 ;
        RECT 72.095 71.905 73.095 72.905 ;
        RECT 77.520 72.370 78.420 72.530 ;
        RECT 77.500 71.730 78.440 72.370 ;
        RECT 77.520 71.570 78.420 71.730 ;
        RECT 49.735 70.990 50.635 71.150 ;
        RECT 49.715 70.350 50.655 70.990 ;
        RECT 49.735 70.190 50.635 70.350 ;
        RECT 56.460 68.405 57.040 69.045 ;
        RECT 56.645 67.700 56.785 68.405 ;
        RECT 72.550 68.235 73.130 68.485 ;
        RECT 73.810 68.235 74.400 68.490 ;
        RECT 61.730 68.020 62.630 68.180 ;
        RECT 72.550 68.095 74.400 68.235 ;
        RECT 56.420 67.050 57.010 67.700 ;
        RECT 61.710 67.380 62.650 68.020 ;
        RECT 72.550 67.845 73.130 68.095 ;
        RECT 73.810 67.840 74.400 68.095 ;
        RECT 61.730 67.220 62.630 67.380 ;
        RECT 49.570 64.885 50.570 65.885 ;
        RECT 49.735 64.450 50.635 64.610 ;
        RECT 49.715 63.810 50.655 64.450 ;
        RECT 49.735 63.650 50.635 63.810 ;
        RECT 56.660 62.365 56.800 67.050 ;
        RECT 61.730 66.200 62.630 66.360 ;
        RECT 61.710 65.560 62.650 66.200 ;
        RECT 74.035 65.975 74.175 67.840 ;
        RECT 61.730 65.400 62.630 65.560 ;
        RECT 73.810 65.325 74.400 65.975 ;
        RECT 61.730 64.380 62.630 64.540 ;
        RECT 61.710 63.740 62.650 64.380 ;
        RECT 61.730 63.580 62.630 63.740 ;
        RECT 74.035 63.370 74.175 65.325 ;
        RECT 61.740 62.565 62.640 62.725 ;
        RECT 73.810 62.720 74.400 63.370 ;
        RECT 56.440 61.715 57.030 62.365 ;
        RECT 61.720 61.925 62.660 62.565 ;
        RECT 61.740 61.765 62.640 61.925 ;
        RECT 46.020 58.780 46.600 59.010 ;
        RECT 43.330 58.640 46.600 58.780 ;
        RECT 28.785 57.165 35.890 57.180 ;
        RECT 28.785 56.525 36.180 57.165 ;
        RECT 28.785 56.480 35.890 56.525 ;
        RECT 28.785 46.505 34.895 56.480 ;
        RECT 28.785 45.805 36.180 46.505 ;
        RECT 28.785 44.950 34.895 45.805 ;
        RECT 35.410 44.950 36.720 45.295 ;
        RECT 28.785 44.250 36.720 44.950 ;
        RECT 41.825 44.525 42.725 44.685 ;
        RECT 28.785 38.370 34.895 44.250 ;
        RECT 35.410 43.925 36.720 44.250 ;
        RECT 41.805 43.885 42.745 44.525 ;
        RECT 41.825 43.725 42.725 43.885 ;
        RECT 43.330 42.150 43.470 58.640 ;
        RECT 46.020 58.370 46.600 58.640 ;
        RECT 49.570 58.195 50.570 59.195 ;
        RECT 49.735 57.755 50.635 57.915 ;
        RECT 49.715 57.115 50.655 57.755 ;
        RECT 49.735 56.955 50.635 57.115 ;
        RECT 56.645 53.880 56.785 61.715 ;
        RECT 61.740 60.740 62.640 60.900 ;
        RECT 74.035 60.840 74.175 62.720 ;
        RECT 61.720 60.100 62.660 60.740 ;
        RECT 73.810 60.190 74.400 60.840 ;
        RECT 61.740 59.940 62.640 60.100 ;
        RECT 61.740 58.915 62.640 59.075 ;
        RECT 61.720 58.275 62.660 58.915 ;
        RECT 61.740 58.115 62.640 58.275 ;
        RECT 74.035 58.195 74.175 60.190 ;
        RECT 73.810 57.545 74.400 58.195 ;
        RECT 61.730 57.105 62.630 57.265 ;
        RECT 61.710 56.465 62.650 57.105 ;
        RECT 61.730 56.305 62.630 56.465 ;
        RECT 74.035 55.720 74.175 57.545 ;
        RECT 59.435 55.280 60.335 55.440 ;
        RECT 61.740 55.280 62.640 55.440 ;
        RECT 59.415 54.640 60.355 55.280 ;
        RECT 61.720 54.640 62.660 55.280 ;
        RECT 73.810 55.070 74.400 55.720 ;
        RECT 71.230 54.795 71.810 55.060 ;
        RECT 72.485 54.795 73.075 55.050 ;
        RECT 71.230 54.655 73.075 54.795 ;
        RECT 59.435 54.480 60.335 54.640 ;
        RECT 61.740 54.480 62.640 54.640 ;
        RECT 71.230 54.420 71.810 54.655 ;
        RECT 72.485 54.400 73.075 54.655 ;
        RECT 84.245 54.325 84.385 75.955 ;
        RECT 109.750 75.700 110.340 76.350 ;
        RECT 113.005 75.920 114.005 76.920 ;
        RECT 114.510 76.545 115.410 76.705 ;
        RECT 114.490 75.905 115.430 76.545 ;
        RECT 114.510 75.745 115.410 75.905 ;
        RECT 93.930 75.540 94.830 75.700 ;
        RECT 92.450 74.440 93.450 75.440 ;
        RECT 93.910 74.900 94.850 75.540 ;
        RECT 112.580 75.295 113.480 75.455 ;
        RECT 93.930 74.740 94.830 74.900 ;
        RECT 111.100 74.195 112.100 75.195 ;
        RECT 112.560 74.655 113.500 75.295 ;
        RECT 112.580 74.495 113.480 74.655 ;
        RECT 91.420 72.875 92.420 73.875 ;
        RECT 92.880 73.870 93.780 74.030 ;
        RECT 92.860 73.230 93.800 73.870 ;
        RECT 92.880 73.070 93.780 73.230 ;
        RECT 110.070 72.630 111.070 73.630 ;
        RECT 111.530 73.625 112.430 73.785 ;
        RECT 111.510 72.985 112.450 73.625 ;
        RECT 111.530 72.825 112.430 72.985 ;
        RECT 87.565 71.475 88.465 71.635 ;
        RECT 87.545 70.835 88.485 71.475 ;
        RECT 89.070 71.370 90.070 72.370 ;
        RECT 90.765 72.290 91.665 72.450 ;
        RECT 90.745 71.650 91.685 72.290 ;
        RECT 90.765 71.490 91.665 71.650 ;
        RECT 106.215 71.230 107.115 71.390 ;
        RECT 87.565 70.675 88.465 70.835 ;
        RECT 106.195 70.590 107.135 71.230 ;
        RECT 107.720 71.125 108.720 72.125 ;
        RECT 109.415 72.045 110.315 72.205 ;
        RECT 109.395 71.405 110.335 72.045 ;
        RECT 109.415 71.245 110.315 71.405 ;
        RECT 106.215 70.430 107.115 70.590 ;
        RECT 85.855 69.230 86.855 70.230 ;
        RECT 87.565 69.115 88.465 69.275 ;
        RECT 87.545 68.475 88.485 69.115 ;
        RECT 104.505 69.000 105.505 70.000 ;
        RECT 124.160 69.870 129.040 87.775 ;
        RECT 120.350 69.170 129.040 69.870 ;
        RECT 106.215 68.870 107.115 69.030 ;
        RECT 87.565 68.315 88.465 68.475 ;
        RECT 106.195 68.230 107.135 68.870 ;
        RECT 106.215 68.070 107.115 68.230 ;
        RECT 88.390 66.830 89.390 67.830 ;
        RECT 89.900 67.650 90.800 67.810 ;
        RECT 89.880 67.010 90.820 67.650 ;
        RECT 89.900 66.850 90.800 67.010 ;
        RECT 107.040 66.585 108.040 67.585 ;
        RECT 108.550 67.405 109.450 67.565 ;
        RECT 108.530 66.765 109.470 67.405 ;
        RECT 108.550 66.605 109.450 66.765 ;
        RECT 90.465 65.405 91.465 66.405 ;
        RECT 92.005 66.130 92.905 66.290 ;
        RECT 91.985 65.490 92.925 66.130 ;
        RECT 92.005 65.330 92.905 65.490 ;
        RECT 109.115 65.160 110.115 66.160 ;
        RECT 110.655 65.885 111.555 66.045 ;
        RECT 110.635 65.245 111.575 65.885 ;
        RECT 110.655 65.085 111.555 65.245 ;
        RECT 90.465 63.460 91.465 64.460 ;
        RECT 92.210 64.305 93.110 64.465 ;
        RECT 92.190 63.665 93.130 64.305 ;
        RECT 102.250 64.115 102.840 64.490 ;
        RECT 92.210 63.505 93.110 63.665 ;
        RECT 92.735 61.920 93.735 62.920 ;
        RECT 94.290 62.845 95.190 63.005 ;
        RECT 94.270 62.205 95.210 62.845 ;
        RECT 94.290 62.045 95.190 62.205 ;
        RECT 95.890 61.920 96.890 62.920 ;
        RECT 102.195 60.025 102.895 64.115 ;
        RECT 109.115 63.215 110.115 64.215 ;
        RECT 110.860 64.060 111.760 64.220 ;
        RECT 110.840 63.420 111.780 64.060 ;
        RECT 110.860 63.260 111.760 63.420 ;
        RECT 111.385 61.675 112.385 62.675 ;
        RECT 112.940 62.600 113.840 62.760 ;
        RECT 112.920 61.960 113.860 62.600 ;
        RECT 112.940 61.800 113.840 61.960 ;
        RECT 114.540 61.675 115.540 62.675 ;
        RECT 124.160 60.025 129.040 69.170 ;
        RECT 102.195 59.325 129.040 60.025 ;
        RECT 102.225 58.655 102.925 59.325 ;
        RECT 73.945 54.185 84.385 54.325 ;
        RECT 99.740 57.955 102.925 58.655 ;
        RECT 56.420 53.230 57.010 53.880 ;
        RECT 73.945 53.845 74.085 54.185 ;
        RECT 58.520 53.705 74.085 53.845 ;
        RECT 49.570 51.530 50.570 52.530 ;
        RECT 49.660 50.825 50.560 50.985 ;
        RECT 49.640 50.185 50.580 50.825 ;
        RECT 49.660 50.025 50.560 50.185 ;
        RECT 56.660 48.310 56.800 53.230 ;
        RECT 58.520 51.695 58.660 53.705 ;
        RECT 99.740 53.060 100.440 57.955 ;
        RECT 105.205 56.970 106.105 57.130 ;
        RECT 105.185 56.330 106.125 56.970 ;
        RECT 105.205 56.170 106.105 56.330 ;
        RECT 106.740 56.040 107.740 57.040 ;
        RECT 108.210 56.970 109.110 57.130 ;
        RECT 108.190 56.330 109.130 56.970 ;
        RECT 108.210 56.170 109.110 56.330 ;
        RECT 109.740 56.040 110.740 57.040 ;
        RECT 112.180 56.970 113.080 57.130 ;
        RECT 112.160 56.330 113.100 56.970 ;
        RECT 112.180 56.170 113.080 56.330 ;
        RECT 104.490 54.630 105.490 55.630 ;
        RECT 69.990 52.360 100.440 53.060 ;
        RECT 104.155 52.955 105.155 53.955 ;
        RECT 105.760 53.895 106.660 54.055 ;
        RECT 105.740 53.255 106.680 53.895 ;
        RECT 105.760 53.095 106.660 53.255 ;
        RECT 58.170 50.685 59.120 51.695 ;
        RECT 61.965 51.315 62.865 51.475 ;
        RECT 58.575 49.135 58.715 50.685 ;
        RECT 61.945 50.675 62.885 51.315 ;
        RECT 71.230 51.015 71.810 51.310 ;
        RECT 72.850 51.015 73.440 51.270 ;
        RECT 71.230 50.875 73.440 51.015 ;
        RECT 59.585 49.640 60.585 50.640 ;
        RECT 61.965 50.515 62.865 50.675 ;
        RECT 71.230 50.670 71.810 50.875 ;
        RECT 72.850 50.620 73.440 50.875 ;
        RECT 73.755 50.870 74.455 52.360 ;
        RECT 104.720 51.720 105.620 51.880 ;
        RECT 104.700 51.080 105.640 51.720 ;
        RECT 104.720 50.920 105.620 51.080 ;
        RECT 73.695 50.590 74.455 50.870 ;
        RECT 73.695 50.450 74.570 50.590 ;
        RECT 124.160 50.580 129.040 59.325 ;
        RECT 73.695 50.170 74.455 50.450 ;
        RECT 61.965 49.495 62.865 49.655 ;
        RECT 58.280 48.495 58.860 49.135 ;
        RECT 61.945 48.855 62.885 49.495 ;
        RECT 56.440 47.660 57.030 48.310 ;
        RECT 59.585 47.755 60.585 48.755 ;
        RECT 61.965 48.695 62.865 48.855 ;
        RECT 71.120 48.755 72.120 49.755 ;
        RECT 73.960 48.280 74.100 50.170 ;
        RECT 104.155 49.335 105.155 50.335 ;
        RECT 119.990 49.880 129.040 50.580 ;
        RECT 104.720 48.440 105.620 48.600 ;
        RECT 61.965 47.675 62.865 47.835 ;
        RECT 61.945 47.035 62.885 47.675 ;
        RECT 73.735 47.630 74.325 48.280 ;
        RECT 104.700 47.800 105.640 48.440 ;
        RECT 104.720 47.640 105.620 47.800 ;
        RECT 59.585 45.930 60.585 46.930 ;
        RECT 61.965 46.875 62.865 47.035 ;
        RECT 71.060 46.185 72.060 47.185 ;
        RECT 49.570 44.905 50.570 45.905 ;
        RECT 61.975 45.855 62.875 46.015 ;
        RECT 61.955 45.215 62.895 45.855 ;
        RECT 73.955 45.725 74.095 47.630 ;
        RECT 61.975 45.055 62.875 45.215 ;
        RECT 73.730 45.075 74.320 45.725 ;
        RECT 104.155 45.585 105.155 46.585 ;
        RECT 105.760 46.400 106.660 46.560 ;
        RECT 105.740 45.760 106.680 46.400 ;
        RECT 105.760 45.600 106.660 45.760 ;
        RECT 46.400 44.520 47.300 44.680 ;
        RECT 46.380 43.880 47.320 44.520 ;
        RECT 59.585 44.055 60.585 45.055 ;
        RECT 61.975 44.035 62.875 44.195 ;
        RECT 46.400 43.720 47.300 43.880 ;
        RECT 61.955 43.395 62.895 44.035 ;
        RECT 71.170 43.680 72.170 44.680 ;
        RECT 61.975 43.235 62.875 43.395 ;
        RECT 44.900 42.380 45.800 42.540 ;
        RECT 43.140 41.500 43.730 42.150 ;
        RECT 44.880 41.740 45.820 42.380 ;
        RECT 59.585 42.235 60.585 43.235 ;
        RECT 73.995 43.160 74.135 45.075 ;
        RECT 104.830 43.980 105.830 44.980 ;
        RECT 105.760 43.270 106.660 43.430 ;
        RECT 73.770 42.510 74.360 43.160 ;
        RECT 105.740 42.630 106.680 43.270 ;
        RECT 61.975 42.210 62.875 42.370 ;
        RECT 44.900 41.580 45.800 41.740 ;
        RECT 37.495 38.675 38.495 39.675 ;
        RECT 35.410 38.370 36.720 38.565 ;
        RECT 28.785 37.670 36.720 38.370 ;
        RECT 41.845 37.865 42.745 38.025 ;
        RECT 28.785 31.875 34.895 37.670 ;
        RECT 35.410 37.195 36.720 37.670 ;
        RECT 41.825 37.225 42.765 37.865 ;
        RECT 41.845 37.065 42.745 37.225 ;
        RECT 43.330 36.075 43.470 41.500 ;
        RECT 53.200 41.085 53.790 41.735 ;
        RECT 61.955 41.570 62.895 42.210 ;
        RECT 46.305 38.685 47.305 39.685 ;
        RECT 46.400 37.890 47.300 38.050 ;
        RECT 46.380 37.250 47.320 37.890 ;
        RECT 46.400 37.090 47.300 37.250 ;
        RECT 53.440 36.075 53.580 41.085 ;
        RECT 59.585 40.495 60.585 41.495 ;
        RECT 61.975 41.410 62.875 41.570 ;
        RECT 71.170 41.070 72.170 42.070 ;
        RECT 73.970 40.600 74.110 42.510 ;
        RECT 105.760 42.470 106.660 42.630 ;
        RECT 107.240 42.490 108.240 43.490 ;
        RECT 108.660 43.245 109.560 43.405 ;
        RECT 108.640 42.605 109.580 43.245 ;
        RECT 108.660 42.445 109.560 42.605 ;
        RECT 109.970 42.530 110.970 43.530 ;
        RECT 112.180 43.500 113.080 43.660 ;
        RECT 112.160 42.860 113.100 43.500 ;
        RECT 124.160 43.480 129.040 49.880 ;
        RECT 123.885 43.430 129.040 43.480 ;
        RECT 112.180 42.700 113.080 42.860 ;
        RECT 123.520 42.790 129.040 43.430 ;
        RECT 123.885 42.780 129.040 42.790 ;
        RECT 61.965 40.400 62.865 40.560 ;
        RECT 61.945 39.760 62.885 40.400 ;
        RECT 73.745 39.950 74.335 40.600 ;
        RECT 110.925 40.440 111.515 41.090 ;
        RECT 59.585 38.660 60.585 39.660 ;
        RECT 61.965 39.600 62.865 39.760 ;
        RECT 61.975 38.575 62.875 38.735 ;
        RECT 71.170 38.585 72.170 39.585 ;
        RECT 61.955 37.935 62.895 38.575 ;
        RECT 61.975 37.775 62.875 37.935 ;
        RECT 71.265 37.550 71.845 37.720 ;
        RECT 68.235 37.250 72.860 37.550 ;
        RECT 43.330 35.930 43.475 36.075 ;
        RECT 53.440 35.930 53.585 36.075 ;
        RECT 43.335 35.445 43.475 35.930 ;
        RECT 43.110 34.795 43.700 35.445 ;
        RECT 44.900 35.415 45.800 35.575 ;
        RECT 35.410 31.875 36.720 32.470 ;
        RECT 37.145 31.970 38.145 32.970 ;
        RECT 28.785 31.175 36.720 31.875 ;
        RECT 41.805 31.750 42.705 31.910 ;
        RECT 21.395 29.645 23.635 29.655 ;
        RECT 28.785 29.645 34.895 31.175 ;
        RECT 35.410 31.100 36.720 31.175 ;
        RECT 41.785 31.110 42.725 31.750 ;
        RECT 41.805 30.950 42.705 31.110 ;
        RECT 21.395 27.645 34.895 29.645 ;
        RECT 43.335 29.355 43.475 34.795 ;
        RECT 44.880 34.775 45.820 35.415 ;
        RECT 53.445 35.400 53.585 35.930 ;
        RECT 55.860 35.825 56.760 35.985 ;
        RECT 44.900 34.615 45.800 34.775 ;
        RECT 53.220 34.750 53.810 35.400 ;
        RECT 55.840 35.185 56.780 35.825 ;
        RECT 55.860 35.025 56.760 35.185 ;
        RECT 46.290 31.980 47.290 32.980 ;
        RECT 47.590 31.730 48.490 31.890 ;
        RECT 47.570 31.090 48.510 31.730 ;
        RECT 47.590 30.930 48.490 31.090 ;
        RECT 53.445 29.375 53.585 34.750 ;
        RECT 57.145 34.450 58.145 35.450 ;
        RECT 64.760 33.690 65.350 33.750 ;
        RECT 64.760 33.100 65.490 33.690 ;
        RECT 57.145 31.405 58.145 32.405 ;
        RECT 43.110 28.705 43.700 29.355 ;
        RECT 44.900 29.130 45.800 29.290 ;
        RECT 21.395 27.455 23.635 27.645 ;
        RECT 28.785 25.650 34.895 27.645 ;
        RECT 35.580 25.650 36.890 26.100 ;
        RECT 37.145 25.855 38.145 26.855 ;
        RECT 28.785 24.950 36.890 25.650 ;
        RECT 41.845 25.325 42.745 25.485 ;
        RECT 28.785 17.065 34.895 24.950 ;
        RECT 35.580 24.730 36.890 24.950 ;
        RECT 41.825 24.685 42.765 25.325 ;
        RECT 41.845 24.525 42.745 24.685 ;
        RECT 43.335 22.880 43.475 28.705 ;
        RECT 44.880 28.490 45.820 29.130 ;
        RECT 53.220 28.725 53.810 29.375 ;
        RECT 44.900 28.330 45.800 28.490 ;
        RECT 46.325 25.885 47.325 26.885 ;
        RECT 47.590 25.325 48.490 25.485 ;
        RECT 47.570 24.685 48.510 25.325 ;
        RECT 47.590 24.525 48.490 24.685 ;
        RECT 44.900 23.055 45.800 23.215 ;
        RECT 43.110 22.230 43.700 22.880 ;
        RECT 44.880 22.415 45.820 23.055 ;
        RECT 53.445 23.030 53.585 28.725 ;
        RECT 55.070 26.415 61.905 27.065 ;
        RECT 44.900 22.255 45.800 22.415 ;
        RECT 53.220 22.380 53.810 23.030 ;
        RECT 36.155 19.460 37.155 20.460 ;
        RECT 43.335 17.995 43.475 22.230 ;
        RECT 46.280 19.480 47.280 20.480 ;
        RECT 53.445 17.995 53.585 22.380 ;
        RECT 43.335 17.855 53.585 17.995 ;
        RECT 55.070 17.065 55.720 26.415 ;
        RECT 61.675 23.995 61.905 25.855 ;
        RECT 61.675 21.575 61.905 23.435 ;
        RECT 28.785 16.415 55.720 17.065 ;
        RECT 28.785 10.600 34.895 16.415 ;
        RECT 64.790 15.865 65.490 33.100 ;
        RECT 68.235 32.200 68.535 37.250 ;
        RECT 71.265 37.080 71.845 37.250 ;
        RECT 72.560 36.340 72.860 37.250 ;
        RECT 73.915 36.920 74.055 39.950 ;
        RECT 111.150 39.610 111.290 40.440 ;
        RECT 110.850 38.970 111.430 39.610 ;
        RECT 74.220 36.920 74.810 37.175 ;
        RECT 73.915 36.780 74.810 36.920 ;
        RECT 74.220 36.525 74.810 36.780 ;
        RECT 71.010 34.805 71.960 35.815 ;
        RECT 72.495 35.700 73.075 36.340 ;
        RECT 68.940 33.910 69.840 34.070 ;
        RECT 68.920 33.270 69.860 33.910 ;
        RECT 68.940 33.110 69.840 33.270 ;
        RECT 71.475 32.200 72.065 32.385 ;
        RECT 68.235 31.900 72.065 32.200 ;
        RECT 71.475 31.735 72.065 31.900 ;
        RECT 55.515 10.585 65.515 15.865 ;
        RECT 78.745 15.680 79.445 33.940 ;
        RECT 86.740 25.205 86.970 27.065 ;
        RECT 86.740 22.785 86.970 24.645 ;
        RECT 86.740 21.575 87.950 22.225 ;
        RECT 87.300 18.435 87.950 21.575 ;
        RECT 95.365 18.435 96.365 18.610 ;
        RECT 87.300 17.785 96.365 18.435 ;
        RECT 87.300 15.850 87.950 17.785 ;
        RECT 95.365 17.610 96.365 17.785 ;
        RECT 124.160 16.840 129.040 42.780 ;
        RECT 138.245 16.840 140.485 16.920 ;
        RECT 69.455 10.605 79.455 15.680 ;
        RECT 86.420 10.610 96.420 15.850 ;
        RECT 124.160 14.840 140.485 16.840 ;
        RECT 63.870 6.215 64.870 10.585 ;
        RECT 77.660 8.120 78.660 10.605 ;
        RECT 91.810 10.060 92.810 10.610 ;
        RECT 124.160 10.600 129.040 14.840 ;
        RECT 138.245 14.720 140.485 14.840 ;
        RECT 138.725 10.060 140.005 10.200 ;
        RECT 91.810 9.060 140.005 10.060 ;
        RECT 138.725 8.960 140.005 9.060 ;
        RECT 77.660 7.990 129.105 8.120 ;
        RECT 77.660 7.120 129.675 7.990 ;
        RECT 128.395 6.750 129.675 7.120 ;
        RECT 63.870 6.070 106.860 6.215 ;
        RECT 63.870 5.215 107.740 6.070 ;
        RECT 106.460 4.830 107.740 5.215 ;
        RECT 14.125 4.405 85.095 4.480 ;
        RECT 14.125 3.855 85.400 4.405 ;
        RECT 14.165 3.480 85.400 3.855 ;
        RECT 84.120 3.165 85.400 3.480 ;
        RECT 9.315 2.865 62.360 3.005 ;
        RECT 9.315 2.005 63.225 2.865 ;
        RECT 61.945 1.625 63.225 2.005 ;
      LAYER met2 ;
        RECT 97.535 212.885 98.265 213.655 ;
        RECT 105.730 213.025 106.460 213.795 ;
        RECT 103.035 210.325 103.615 210.425 ;
        RECT 106.955 210.325 107.535 210.425 ;
        RECT 64.085 210.045 64.665 210.215 ;
        RECT 93.170 210.045 93.750 210.215 ;
        RECT 103.035 210.185 107.535 210.325 ;
        RECT 64.085 209.745 95.280 210.045 ;
        RECT 103.035 209.785 103.615 210.185 ;
        RECT 64.085 209.575 64.665 209.745 ;
        RECT 93.170 209.575 93.750 209.745 ;
        RECT 53.510 209.085 54.090 209.285 ;
        RECT 53.510 208.785 60.815 209.085 ;
        RECT 53.510 208.645 54.090 208.785 ;
        RECT 53.470 204.245 54.050 204.475 ;
        RECT 60.515 204.245 60.815 208.785 ;
        RECT 63.905 206.260 64.485 206.410 ;
        RECT 93.170 206.260 93.750 206.430 ;
        RECT 63.905 205.960 93.750 206.260 ;
        RECT 63.905 205.770 64.485 205.960 ;
        RECT 93.170 205.790 93.750 205.960 ;
        RECT 64.045 205.295 64.345 205.770 ;
        RECT 63.905 204.655 64.485 205.295 ;
        RECT 53.470 203.945 76.620 204.245 ;
        RECT 53.470 203.835 54.050 203.945 ;
        RECT 76.320 201.005 76.620 203.945 ;
        RECT 76.220 200.365 76.800 201.005 ;
        RECT 53.180 189.405 54.310 190.575 ;
        RECT 56.630 186.520 57.210 187.160 ;
        RECT 54.445 184.640 55.025 184.810 ;
        RECT 56.775 184.640 57.075 186.520 ;
        RECT 54.445 184.340 57.075 184.640 ;
        RECT 54.445 184.170 55.025 184.340 ;
        RECT 89.235 176.030 89.815 176.200 ;
        RECT 89.235 175.990 93.535 176.030 ;
        RECT 94.980 175.990 95.280 209.745 ;
        RECT 97.535 205.710 98.265 206.480 ;
        RECT 103.120 203.110 103.700 203.360 ;
        RECT 105.265 203.110 105.405 210.185 ;
        RECT 106.955 209.785 107.535 210.185 ;
        RECT 105.730 205.945 106.460 206.715 ;
        RECT 107.040 203.110 107.620 203.360 ;
        RECT 103.120 202.970 107.620 203.110 ;
        RECT 103.120 202.720 103.700 202.970 ;
        RECT 97.535 198.760 98.265 199.530 ;
        RECT 103.120 196.230 103.700 196.480 ;
        RECT 105.265 196.230 105.405 202.970 ;
        RECT 107.040 202.720 107.620 202.970 ;
        RECT 105.730 199.075 106.460 199.845 ;
        RECT 107.040 196.230 107.620 196.480 ;
        RECT 103.120 196.090 107.620 196.230 ;
        RECT 103.120 195.840 103.700 196.090 ;
        RECT 95.765 191.685 96.495 192.455 ;
        RECT 97.535 191.735 98.265 192.505 ;
        RECT 97.535 189.070 98.265 189.475 ;
        RECT 103.120 189.070 103.700 189.320 ;
        RECT 105.265 189.070 105.405 196.090 ;
        RECT 107.040 195.840 107.620 196.090 ;
        RECT 105.730 191.735 106.460 192.505 ;
        RECT 107.040 189.070 107.620 189.320 ;
        RECT 97.535 188.930 107.620 189.070 ;
        RECT 97.535 188.705 98.265 188.930 ;
        RECT 103.120 188.680 103.700 188.930 ;
        RECT 107.040 188.680 107.620 188.930 ;
        RECT 89.235 175.730 95.280 175.990 ;
        RECT 89.235 175.560 89.815 175.730 ;
        RECT 93.235 175.690 95.280 175.730 ;
        RECT 89.260 172.015 89.840 172.230 ;
        RECT 86.220 171.715 89.840 172.015 ;
        RECT 52.745 170.140 53.445 170.145 ;
        RECT 52.515 169.440 55.235 170.140 ;
        RECT 52.535 165.460 53.115 165.465 ;
        RECT 54.535 165.460 55.235 169.440 ;
        RECT 52.535 164.825 55.235 165.460 ;
        RECT 52.575 164.760 55.235 164.825 ;
        RECT 52.540 160.700 53.435 160.715 ;
        RECT 54.535 160.700 55.235 164.760 ;
        RECT 86.220 162.085 86.520 171.715 ;
        RECT 89.260 171.590 89.840 171.715 ;
        RECT 89.250 165.970 89.830 166.140 ;
        RECT 93.235 165.970 93.535 175.690 ;
        RECT 105.700 172.670 106.430 173.440 ;
        RECT 93.975 165.970 94.555 166.170 ;
        RECT 89.250 165.670 94.555 165.970 ;
        RECT 105.700 165.880 106.430 166.650 ;
        RECT 89.250 165.500 89.830 165.670 ;
        RECT 93.975 165.530 94.555 165.670 ;
        RECT 86.115 162.070 86.695 162.085 ;
        RECT 89.260 162.070 89.840 162.240 ;
        RECT 86.115 161.770 89.840 162.070 ;
        RECT 86.115 161.445 86.695 161.770 ;
        RECT 89.260 161.600 89.840 161.770 ;
        RECT 55.415 160.700 56.115 160.715 ;
        RECT 52.480 160.000 56.115 160.700 ;
        RECT 21.330 146.470 23.700 148.800 ;
        RECT 138.180 145.485 140.550 147.815 ;
        RECT 52.155 109.025 81.015 109.165 ;
        RECT 44.050 108.110 44.950 108.300 ;
        RECT 41.595 107.410 44.950 108.110 ;
        RECT 41.595 105.785 42.295 107.410 ;
        RECT 44.050 107.340 44.950 107.410 ;
        RECT 52.155 107.900 52.295 109.025 ;
        RECT 53.035 107.900 53.935 108.310 ;
        RECT 52.155 107.760 53.935 107.900 ;
        RECT 41.595 104.825 43.195 105.785 ;
        RECT 41.595 99.435 42.295 104.825 ;
        RECT 43.910 101.070 45.040 102.240 ;
        RECT 44.050 99.435 44.950 99.450 ;
        RECT 41.595 98.735 44.950 99.435 ;
        RECT 41.595 95.990 42.295 98.735 ;
        RECT 43.920 98.700 44.950 98.735 ;
        RECT 44.050 98.490 44.950 98.700 ;
        RECT 52.155 97.850 52.295 107.760 ;
        RECT 53.035 107.350 53.935 107.760 ;
        RECT 62.340 107.900 62.480 109.025 ;
        RECT 63.270 107.900 64.170 108.310 ;
        RECT 71.600 108.060 72.330 108.830 ;
        RECT 76.775 108.775 77.675 108.835 ;
        RECT 76.775 108.075 79.730 108.775 ;
        RECT 62.340 107.760 64.170 107.900 ;
        RECT 76.775 107.875 77.675 108.075 ;
        RECT 59.510 105.510 60.410 105.640 ;
        RECT 59.490 104.680 60.410 105.510 ;
        RECT 52.895 101.105 54.025 102.275 ;
        RECT 53.035 97.850 53.935 98.350 ;
        RECT 52.145 97.710 53.935 97.850 ;
        RECT 41.595 95.030 43.195 95.990 ;
        RECT 35.375 88.415 35.955 88.425 ;
        RECT 41.595 88.415 42.295 95.030 ;
        RECT 43.910 91.160 45.040 92.330 ;
        RECT 35.375 88.230 44.500 88.415 ;
        RECT 35.375 87.785 44.950 88.230 ;
        RECT 52.155 88.170 52.295 97.710 ;
        RECT 53.035 97.390 53.935 97.710 ;
        RECT 59.490 95.290 60.190 104.680 ;
        RECT 62.340 97.870 62.480 107.760 ;
        RECT 63.270 107.350 64.170 107.760 ;
        RECT 79.030 106.820 79.730 108.075 ;
        RECT 79.030 106.120 80.600 106.820 ;
        RECT 69.535 104.680 70.435 105.640 ;
        RECT 63.390 101.045 64.520 102.215 ;
        RECT 63.270 97.870 64.170 98.370 ;
        RECT 62.340 97.730 64.170 97.870 ;
        RECT 59.490 94.330 60.410 95.290 ;
        RECT 52.895 91.195 54.025 92.365 ;
        RECT 53.035 88.170 53.935 88.580 ;
        RECT 52.145 88.030 53.935 88.170 ;
        RECT 35.665 87.715 44.950 87.785 ;
        RECT 41.595 86.630 42.295 87.715 ;
        RECT 44.050 87.270 44.950 87.715 ;
        RECT 41.595 85.670 43.195 86.630 ;
        RECT 41.595 78.985 42.295 85.670 ;
        RECT 43.910 81.005 45.040 82.175 ;
        RECT 44.050 78.985 44.950 79.155 ;
        RECT 41.595 78.285 44.950 78.985 ;
        RECT 52.155 78.705 52.295 88.030 ;
        RECT 53.035 87.620 53.935 88.030 ;
        RECT 59.490 85.270 60.190 94.330 ;
        RECT 62.340 88.295 62.480 97.730 ;
        RECT 63.270 97.410 64.170 97.730 ;
        RECT 69.635 95.290 70.335 104.680 ;
        RECT 77.425 101.795 78.325 101.925 ;
        RECT 77.410 100.965 78.325 101.795 ;
        RECT 77.410 100.825 78.110 100.965 ;
        RECT 79.030 100.825 79.730 106.120 ;
        RECT 79.900 106.105 80.600 106.120 ;
        RECT 80.875 105.050 81.015 109.025 ;
        RECT 80.365 104.660 81.015 105.050 ;
        RECT 80.365 104.410 80.945 104.660 ;
        RECT 76.770 100.125 79.730 100.825 ;
        RECT 76.770 98.835 77.470 100.125 ;
        RECT 76.700 97.875 77.600 98.835 ;
        RECT 69.535 94.330 70.435 95.290 ;
        RECT 63.390 91.150 64.520 92.320 ;
        RECT 63.270 88.295 64.170 88.705 ;
        RECT 62.340 88.155 64.170 88.295 ;
        RECT 59.490 84.310 60.410 85.270 ;
        RECT 52.895 81.180 54.025 82.350 ;
        RECT 53.035 78.705 53.935 79.145 ;
        RECT 52.155 78.565 53.935 78.705 ;
        RECT 41.595 76.145 42.295 78.285 ;
        RECT 44.050 78.195 44.950 78.285 ;
        RECT 53.035 78.185 53.935 78.565 ;
        RECT 59.490 76.335 60.190 84.310 ;
        RECT 62.340 78.735 62.480 88.155 ;
        RECT 63.270 87.745 64.170 88.155 ;
        RECT 69.635 85.430 70.335 94.330 ;
        RECT 77.425 91.445 78.325 92.405 ;
        RECT 77.525 90.550 78.225 91.445 ;
        RECT 79.030 90.550 79.730 100.125 ;
        RECT 120.135 97.140 120.865 97.910 ;
        RECT 94.125 96.000 114.980 96.140 ;
        RECT 94.125 93.990 94.265 96.000 ;
        RECT 94.580 94.370 95.710 95.540 ;
        RECT 96.470 95.240 96.610 96.000 ;
        RECT 96.150 94.280 97.050 95.240 ;
        RECT 92.675 92.645 93.805 93.815 ;
        RECT 94.125 93.440 95.120 93.990 ;
        RECT 94.220 93.030 95.120 93.440 ;
        RECT 76.745 89.850 79.730 90.550 ;
        RECT 88.235 91.425 91.150 91.565 ;
        RECT 88.235 89.925 88.375 91.425 ;
        RECT 76.745 89.005 77.445 89.850 ;
        RECT 76.700 88.045 77.600 89.005 ;
        RECT 69.535 84.470 70.435 85.430 ;
        RECT 63.390 81.295 64.520 82.465 ;
        RECT 63.270 78.735 64.170 79.190 ;
        RECT 62.340 78.595 64.170 78.735 ;
        RECT 63.270 78.230 64.170 78.595 ;
        RECT 41.595 75.315 42.590 76.145 ;
        RECT 41.690 75.185 42.590 75.315 ;
        RECT 50.465 75.235 51.195 76.005 ;
        RECT 59.490 75.375 60.410 76.335 ;
        RECT 69.635 76.105 70.335 84.470 ;
        RECT 72.435 81.445 73.565 82.615 ;
        RECT 77.390 81.090 78.290 82.050 ;
        RECT 77.565 80.355 78.265 81.090 ;
        RECT 79.030 80.355 79.730 89.850 ;
        RECT 87.855 88.965 88.755 89.925 ;
        RECT 89.295 89.575 90.425 90.745 ;
        RECT 91.010 90.740 91.150 91.425 ;
        RECT 91.645 91.080 92.775 92.250 ;
        RECT 93.170 91.910 94.070 92.320 ;
        RECT 94.510 91.910 94.650 93.030 ;
        RECT 93.170 91.770 94.650 91.910 ;
        RECT 93.170 91.360 94.070 91.770 ;
        RECT 91.010 90.525 91.955 90.740 ;
        RECT 93.550 90.525 93.690 91.360 ;
        RECT 91.010 90.385 93.690 90.525 ;
        RECT 91.010 90.190 91.955 90.385 ;
        RECT 91.055 89.780 91.955 90.190 ;
        RECT 86.080 87.415 87.210 88.585 ;
        RECT 88.235 87.565 88.375 88.965 ;
        RECT 87.855 87.155 88.755 87.565 ;
        RECT 87.815 86.605 88.755 87.155 ;
        RECT 87.815 84.375 87.955 86.605 ;
        RECT 88.615 85.035 89.745 86.205 ;
        RECT 90.190 85.655 91.090 86.100 ;
        RECT 90.190 85.515 92.815 85.655 ;
        RECT 90.190 85.140 91.090 85.515 ;
        RECT 90.335 84.375 90.475 85.140 ;
        RECT 87.815 84.235 90.475 84.375 ;
        RECT 89.830 81.095 89.970 84.235 ;
        RECT 90.690 83.610 91.820 84.780 ;
        RECT 92.675 84.580 92.815 85.515 ;
        RECT 92.295 83.620 93.195 84.580 ;
        RECT 90.690 81.665 91.820 82.835 ;
        RECT 92.500 82.345 93.400 82.755 ;
        RECT 92.415 81.795 93.400 82.345 ;
        RECT 92.415 81.095 92.555 81.795 ;
        RECT 89.830 80.955 92.555 81.095 ;
        RECT 76.930 79.655 79.730 80.355 ;
        RECT 76.930 78.880 77.630 79.655 ;
        RECT 76.860 77.920 77.760 78.880 ;
        RECT 43.910 72.000 45.040 73.170 ;
        RECT 52.895 71.975 54.025 73.145 ;
        RECT 49.735 71.130 50.635 71.150 ;
        RECT 49.005 70.990 50.635 71.130 ;
        RECT 49.005 64.565 49.145 70.990 ;
        RECT 49.735 70.190 50.635 70.990 ;
        RECT 59.490 70.140 60.190 75.375 ;
        RECT 69.535 75.145 70.435 76.105 ;
        RECT 63.390 72.120 64.520 73.290 ;
        RECT 69.635 70.140 70.335 75.145 ;
        RECT 72.030 71.820 73.160 72.990 ;
        RECT 77.520 71.570 78.420 72.530 ;
        RECT 77.685 70.140 78.385 71.570 ;
        RECT 79.030 70.140 79.730 79.655 ;
        RECT 91.480 79.355 91.620 80.955 ;
        RECT 92.960 80.125 94.090 81.295 ;
        RECT 94.580 80.335 95.480 81.295 ;
        RECT 94.960 79.355 95.100 80.335 ;
        RECT 96.115 80.125 97.245 81.295 ;
        RECT 91.480 79.215 95.100 79.355 ;
        RECT 102.225 77.605 102.365 96.000 ;
        RECT 112.455 93.990 112.595 96.000 ;
        RECT 112.910 94.370 114.040 95.540 ;
        RECT 114.840 95.240 114.980 96.000 ;
        RECT 114.480 94.280 115.380 95.240 ;
        RECT 102.710 91.960 103.840 93.130 ;
        RECT 111.005 92.645 112.135 93.815 ;
        RECT 112.455 93.440 113.450 93.990 ;
        RECT 112.550 93.030 113.450 93.440 ;
        RECT 106.565 91.425 109.480 91.565 ;
        RECT 106.565 89.925 106.705 91.425 ;
        RECT 106.185 88.965 107.085 89.925 ;
        RECT 107.625 89.575 108.755 90.745 ;
        RECT 109.340 90.740 109.480 91.425 ;
        RECT 109.975 91.080 111.105 92.250 ;
        RECT 111.500 91.910 112.400 92.320 ;
        RECT 112.840 91.910 112.980 93.030 ;
        RECT 111.500 91.770 112.980 91.910 ;
        RECT 111.500 91.360 112.400 91.770 ;
        RECT 109.340 90.525 110.285 90.740 ;
        RECT 111.880 90.525 112.020 91.360 ;
        RECT 109.340 90.385 112.020 90.525 ;
        RECT 109.340 90.190 110.285 90.385 ;
        RECT 109.385 89.780 110.285 90.190 ;
        RECT 104.410 87.435 105.540 88.605 ;
        RECT 106.565 87.565 106.705 88.965 ;
        RECT 106.185 87.155 107.085 87.565 ;
        RECT 106.145 86.605 107.085 87.155 ;
        RECT 106.145 84.375 106.285 86.605 ;
        RECT 106.945 85.035 108.075 86.205 ;
        RECT 108.520 85.655 109.420 86.100 ;
        RECT 108.520 85.515 111.145 85.655 ;
        RECT 108.520 85.140 109.420 85.515 ;
        RECT 108.665 84.375 108.805 85.140 ;
        RECT 106.145 84.235 108.805 84.375 ;
        RECT 108.160 81.095 108.300 84.235 ;
        RECT 109.020 83.610 110.150 84.780 ;
        RECT 111.005 84.580 111.145 85.515 ;
        RECT 110.625 83.620 111.525 84.580 ;
        RECT 109.020 81.665 110.150 82.835 ;
        RECT 110.830 82.345 111.730 82.755 ;
        RECT 110.745 81.795 111.730 82.345 ;
        RECT 110.745 81.095 110.885 81.795 ;
        RECT 108.160 80.955 110.885 81.095 ;
        RECT 109.810 79.355 109.950 80.955 ;
        RECT 111.290 80.125 112.420 81.295 ;
        RECT 112.910 80.335 113.810 81.295 ;
        RECT 113.290 79.355 113.430 80.335 ;
        RECT 114.445 80.125 115.575 81.295 ;
        RECT 109.810 79.215 113.430 79.355 ;
        RECT 94.050 77.465 114.970 77.605 ;
        RECT 94.050 75.700 94.190 77.465 ;
        RECT 94.340 76.080 95.470 77.250 ;
        RECT 96.065 76.950 96.205 77.465 ;
        RECT 95.860 75.990 96.760 76.950 ;
        RECT 92.385 74.355 93.515 75.525 ;
        RECT 93.930 74.740 94.830 75.700 ;
        RECT 112.485 75.455 112.625 77.465 ;
        RECT 112.940 75.835 114.070 77.005 ;
        RECT 114.830 76.705 114.970 77.465 ;
        RECT 114.510 75.745 115.410 76.705 ;
        RECT 87.945 73.135 90.860 73.275 ;
        RECT 87.945 71.635 88.085 73.135 ;
        RECT 87.565 70.675 88.465 71.635 ;
        RECT 89.005 71.285 90.135 72.455 ;
        RECT 90.720 72.450 90.860 73.135 ;
        RECT 91.355 72.790 92.485 73.960 ;
        RECT 92.880 73.620 93.780 74.030 ;
        RECT 94.220 73.620 94.360 74.740 ;
        RECT 111.035 74.110 112.165 75.280 ;
        RECT 112.485 74.905 113.480 75.455 ;
        RECT 112.580 74.495 113.480 74.905 ;
        RECT 92.880 73.480 94.360 73.620 ;
        RECT 92.880 73.070 93.780 73.480 ;
        RECT 90.720 72.235 91.665 72.450 ;
        RECT 93.260 72.235 93.400 73.070 ;
        RECT 90.720 72.095 93.400 72.235 ;
        RECT 106.595 72.890 109.510 73.030 ;
        RECT 90.720 71.900 91.665 72.095 ;
        RECT 90.765 71.490 91.665 71.900 ;
        RECT 106.595 71.390 106.735 72.890 ;
        RECT 59.490 69.440 79.730 70.140 ;
        RECT 56.385 68.340 57.115 69.110 ;
        RECT 61.115 67.770 61.255 69.440 ;
        RECT 61.730 67.770 62.630 68.180 ;
        RECT 72.490 67.845 73.190 69.440 ;
        RECT 85.790 69.145 86.920 70.315 ;
        RECT 87.945 69.275 88.085 70.675 ;
        RECT 106.215 70.430 107.115 71.390 ;
        RECT 107.655 71.040 108.785 72.210 ;
        RECT 109.370 72.205 109.510 72.890 ;
        RECT 110.005 72.545 111.135 73.715 ;
        RECT 111.530 73.375 112.430 73.785 ;
        RECT 112.870 73.375 113.010 74.495 ;
        RECT 111.530 73.235 113.010 73.375 ;
        RECT 111.530 72.825 112.430 73.235 ;
        RECT 109.370 71.990 110.315 72.205 ;
        RECT 111.910 71.990 112.050 72.825 ;
        RECT 109.370 71.850 112.050 71.990 ;
        RECT 109.370 71.655 110.315 71.850 ;
        RECT 109.415 71.245 110.315 71.655 ;
        RECT 87.565 68.865 88.465 69.275 ;
        RECT 104.440 68.915 105.570 70.085 ;
        RECT 106.595 69.030 106.735 70.430 ;
        RECT 87.525 68.315 88.465 68.865 ;
        RECT 106.215 68.620 107.115 69.030 ;
        RECT 61.115 67.630 62.630 67.770 ;
        RECT 49.505 64.800 50.635 65.970 ;
        RECT 61.115 65.800 61.255 67.630 ;
        RECT 61.730 67.220 62.630 67.630 ;
        RECT 61.730 65.800 62.630 66.360 ;
        RECT 61.115 65.660 62.630 65.800 ;
        RECT 87.525 65.710 87.665 68.315 ;
        RECT 106.175 68.070 107.115 68.620 ;
        RECT 88.325 66.745 89.455 67.915 ;
        RECT 89.900 66.990 90.800 67.810 ;
        RECT 89.900 66.850 92.525 66.990 ;
        RECT 90.045 65.710 90.185 66.850 ;
        RECT 49.735 64.565 50.635 64.610 ;
        RECT 49.005 64.425 50.635 64.565 ;
        RECT 45.945 58.305 46.675 59.075 ;
        RECT 49.005 57.845 49.145 64.425 ;
        RECT 49.735 63.650 50.635 64.425 ;
        RECT 61.115 64.150 61.255 65.660 ;
        RECT 61.730 65.400 62.630 65.660 ;
        RECT 83.450 65.570 90.185 65.710 ;
        RECT 61.730 64.150 62.630 64.540 ;
        RECT 61.115 64.010 62.630 64.150 ;
        RECT 61.115 62.285 61.255 64.010 ;
        RECT 61.730 63.580 62.630 64.010 ;
        RECT 61.740 62.285 62.640 62.725 ;
        RECT 61.115 62.145 62.640 62.285 ;
        RECT 61.115 60.480 61.255 62.145 ;
        RECT 61.740 61.765 62.640 62.145 ;
        RECT 61.740 60.480 62.640 60.900 ;
        RECT 61.115 60.340 62.640 60.480 ;
        RECT 49.505 58.110 50.635 59.280 ;
        RECT 61.115 58.655 61.255 60.340 ;
        RECT 61.740 59.940 62.640 60.340 ;
        RECT 61.740 58.655 62.640 59.075 ;
        RECT 61.115 58.515 62.640 58.655 ;
        RECT 49.735 57.845 50.635 57.915 ;
        RECT 49.005 57.705 50.635 57.845 ;
        RECT 49.005 57.195 49.145 57.705 ;
        RECT 35.600 56.495 49.145 57.195 ;
        RECT 49.735 56.955 50.635 57.705 ;
        RECT 49.005 50.955 49.145 56.495 ;
        RECT 61.115 56.730 61.255 58.515 ;
        RECT 61.740 58.115 62.640 58.515 ;
        RECT 61.730 56.730 62.630 57.265 ;
        RECT 61.115 56.590 62.630 56.730 ;
        RECT 59.435 54.480 60.335 55.440 ;
        RECT 61.115 55.105 61.255 56.590 ;
        RECT 61.730 56.305 62.630 56.590 ;
        RECT 61.740 55.105 62.640 55.440 ;
        RECT 61.115 54.965 62.640 55.105 ;
        RECT 61.740 54.480 62.640 54.965 ;
        RECT 59.815 52.970 59.955 54.480 ;
        RECT 71.155 54.355 71.885 55.125 ;
        RECT 59.815 52.830 62.465 52.970 ;
        RECT 49.505 51.445 50.635 52.615 ;
        RECT 62.325 51.475 62.465 52.830 ;
        RECT 61.965 51.075 62.865 51.475 ;
        RECT 49.660 50.955 50.560 50.985 ;
        RECT 49.005 50.815 50.560 50.955 ;
        RECT 49.660 50.025 50.560 50.815 ;
        RECT 61.350 50.935 62.865 51.075 ;
        RECT 59.520 49.555 60.650 50.725 ;
        RECT 58.005 48.230 59.135 49.400 ;
        RECT 61.350 49.095 61.490 50.935 ;
        RECT 61.965 50.515 62.865 50.935 ;
        RECT 71.155 50.605 71.885 51.375 ;
        RECT 61.965 49.095 62.865 49.655 ;
        RECT 61.350 48.955 62.865 49.095 ;
        RECT 59.520 47.670 60.650 48.840 ;
        RECT 61.350 47.445 61.490 48.955 ;
        RECT 61.965 48.695 62.865 48.955 ;
        RECT 71.055 48.670 72.185 49.840 ;
        RECT 61.965 47.445 62.865 47.835 ;
        RECT 61.350 47.305 62.865 47.445 ;
        RECT 35.540 46.425 36.240 46.475 ;
        RECT 35.540 45.725 42.625 46.425 ;
        RECT 41.925 44.685 42.625 45.725 ;
        RECT 49.505 44.820 50.635 45.990 ;
        RECT 59.520 45.845 60.650 47.015 ;
        RECT 61.350 45.580 61.490 47.305 ;
        RECT 61.965 46.875 62.865 47.305 ;
        RECT 70.995 46.100 72.125 47.270 ;
        RECT 61.975 45.580 62.875 46.015 ;
        RECT 61.350 45.440 62.875 45.580 ;
        RECT 41.825 44.550 42.725 44.685 ;
        RECT 46.400 44.565 47.300 44.680 ;
        RECT 46.400 44.550 54.855 44.565 ;
        RECT 41.825 43.865 54.855 44.550 ;
        RECT 59.520 43.970 60.650 45.140 ;
        RECT 41.825 43.850 47.300 43.865 ;
        RECT 41.825 43.725 42.725 43.850 ;
        RECT 37.430 38.590 38.560 39.760 ;
        RECT 41.845 37.695 42.745 38.025 ;
        RECT 42.955 37.695 43.095 43.850 ;
        RECT 41.845 37.395 43.095 37.695 ;
        RECT 41.845 37.065 42.745 37.395 ;
        RECT 37.080 31.885 38.210 33.055 ;
        RECT 41.805 31.375 42.705 31.910 ;
        RECT 42.955 31.375 43.095 37.395 ;
        RECT 41.805 31.075 43.095 31.375 ;
        RECT 41.805 30.950 42.705 31.075 ;
        RECT 21.330 27.390 23.700 29.720 ;
        RECT 37.080 25.770 38.210 26.940 ;
        RECT 41.845 24.885 42.745 25.485 ;
        RECT 42.955 24.885 43.095 31.075 ;
        RECT 41.845 24.745 43.095 24.885 ;
        RECT 44.400 42.210 44.700 43.850 ;
        RECT 46.400 43.720 47.300 43.850 ;
        RECT 44.900 42.210 45.800 42.540 ;
        RECT 44.400 41.910 45.800 42.210 ;
        RECT 44.400 37.720 44.700 41.910 ;
        RECT 44.900 41.580 45.800 41.910 ;
        RECT 46.240 38.600 47.370 39.770 ;
        RECT 46.400 37.720 47.300 38.050 ;
        RECT 44.400 37.420 47.300 37.720 ;
        RECT 44.400 35.245 44.700 37.420 ;
        RECT 46.400 37.090 47.300 37.420 ;
        RECT 54.155 35.855 54.855 43.865 ;
        RECT 61.350 43.775 61.490 45.440 ;
        RECT 61.975 45.055 62.875 45.440 ;
        RECT 61.975 43.775 62.875 44.195 ;
        RECT 61.350 43.635 62.875 43.775 ;
        RECT 59.520 42.150 60.650 43.320 ;
        RECT 61.350 41.950 61.490 43.635 ;
        RECT 61.975 43.235 62.875 43.635 ;
        RECT 71.105 43.595 72.235 44.765 ;
        RECT 61.975 41.950 62.875 42.370 ;
        RECT 61.350 41.810 62.875 41.950 ;
        RECT 59.520 40.410 60.650 41.580 ;
        RECT 61.350 40.145 61.490 41.810 ;
        RECT 61.975 41.410 62.875 41.810 ;
        RECT 71.105 40.985 72.235 42.155 ;
        RECT 61.965 40.145 62.865 40.560 ;
        RECT 61.350 40.005 62.865 40.145 ;
        RECT 59.520 38.575 60.650 39.745 ;
        RECT 61.350 38.325 61.490 40.005 ;
        RECT 61.965 39.600 62.865 40.005 ;
        RECT 61.975 38.325 62.875 38.735 ;
        RECT 71.105 38.500 72.235 39.670 ;
        RECT 61.350 38.185 62.875 38.325 ;
        RECT 61.975 37.775 62.875 38.185 ;
        RECT 71.190 37.015 71.920 37.785 ;
        RECT 83.450 37.265 83.590 65.570 ;
        RECT 89.710 62.855 89.850 65.570 ;
        RECT 90.400 65.320 91.530 66.490 ;
        RECT 92.385 66.290 92.525 66.850 ;
        RECT 92.005 65.330 92.905 66.290 ;
        RECT 106.175 65.840 106.315 68.070 ;
        RECT 106.975 66.500 108.105 67.670 ;
        RECT 108.550 67.120 109.450 67.565 ;
        RECT 108.550 66.980 111.175 67.120 ;
        RECT 108.550 66.605 109.450 66.980 ;
        RECT 108.695 65.840 108.835 66.605 ;
        RECT 106.175 65.700 108.835 65.840 ;
        RECT 90.400 63.375 91.530 64.545 ;
        RECT 92.210 64.055 93.110 64.465 ;
        RECT 91.920 63.915 93.110 64.055 ;
        RECT 91.920 62.855 92.060 63.915 ;
        RECT 92.210 63.505 93.110 63.915 ;
        RECT 89.710 62.715 92.060 62.855 ;
        RECT 91.190 60.690 91.330 62.715 ;
        RECT 92.670 61.835 93.800 63.005 ;
        RECT 94.290 62.045 95.190 63.005 ;
        RECT 94.670 60.690 94.810 62.045 ;
        RECT 95.825 61.835 96.955 63.005 ;
        RECT 108.190 62.560 108.330 65.700 ;
        RECT 109.050 65.075 110.180 66.245 ;
        RECT 111.035 66.045 111.175 66.980 ;
        RECT 110.655 65.085 111.555 66.045 ;
        RECT 109.050 63.130 110.180 64.300 ;
        RECT 110.860 63.810 111.760 64.220 ;
        RECT 110.775 63.260 111.760 63.810 ;
        RECT 110.775 62.560 110.915 63.260 ;
        RECT 108.190 62.420 110.915 62.560 ;
        RECT 91.190 60.550 94.810 60.690 ;
        RECT 109.840 60.820 109.980 62.420 ;
        RECT 111.320 61.590 112.450 62.760 ;
        RECT 112.940 61.800 113.840 62.760 ;
        RECT 113.320 60.820 113.460 61.800 ;
        RECT 114.475 61.590 115.605 62.760 ;
        RECT 109.840 60.680 113.460 60.820 ;
        RECT 94.670 60.455 94.810 60.550 ;
        RECT 94.670 60.315 94.850 60.455 ;
        RECT 94.710 59.400 94.850 60.315 ;
        RECT 94.710 59.260 101.790 59.400 ;
        RECT 101.650 39.360 101.790 59.260 ;
        RECT 105.305 57.660 112.980 58.360 ;
        RECT 105.305 57.130 106.005 57.660 ;
        RECT 108.335 57.130 109.035 57.660 ;
        RECT 112.280 57.130 112.980 57.660 ;
        RECT 105.205 57.000 106.105 57.130 ;
        RECT 102.775 56.300 106.105 57.000 ;
        RECT 102.775 51.750 103.475 56.300 ;
        RECT 105.205 56.170 106.105 56.300 ;
        RECT 106.675 55.955 107.805 57.125 ;
        RECT 108.210 56.170 109.110 57.130 ;
        RECT 109.675 55.955 110.805 57.125 ;
        RECT 112.180 56.170 113.080 57.130 ;
        RECT 104.425 54.545 105.555 55.715 ;
        RECT 104.090 52.870 105.220 54.040 ;
        RECT 105.760 53.095 106.660 54.055 ;
        RECT 105.960 52.075 106.660 53.095 ;
        RECT 104.820 51.880 106.660 52.075 ;
        RECT 104.720 51.750 106.660 51.880 ;
        RECT 102.715 51.375 106.660 51.750 ;
        RECT 102.715 51.050 105.620 51.375 ;
        RECT 102.715 48.470 103.415 51.050 ;
        RECT 104.720 50.920 105.620 51.050 ;
        RECT 104.090 49.250 105.220 50.420 ;
        RECT 104.720 48.470 105.620 48.600 ;
        RECT 102.715 48.265 105.620 48.470 ;
        RECT 102.700 47.770 105.620 48.265 ;
        RECT 102.700 47.565 103.415 47.770 ;
        RECT 104.720 47.640 105.620 47.770 ;
        RECT 102.700 41.940 103.400 47.565 ;
        RECT 104.090 45.500 105.220 46.670 ;
        RECT 105.760 45.600 106.660 46.560 ;
        RECT 104.765 43.895 105.895 45.065 ;
        RECT 106.140 43.430 106.280 45.600 ;
        RECT 105.760 42.470 106.660 43.430 ;
        RECT 106.125 41.940 106.265 42.470 ;
        RECT 107.175 42.405 108.305 43.575 ;
        RECT 108.660 42.445 109.560 43.405 ;
        RECT 109.905 42.445 111.035 43.615 ;
        RECT 112.180 43.480 113.080 43.660 ;
        RECT 112.180 43.430 123.885 43.480 ;
        RECT 112.180 42.790 124.110 43.430 ;
        RECT 112.180 42.780 123.885 42.790 ;
        RECT 112.180 42.700 113.080 42.780 ;
        RECT 102.700 41.695 106.615 41.940 ;
        RECT 108.725 41.695 109.425 42.445 ;
        RECT 112.280 41.695 112.980 42.700 ;
        RECT 102.700 41.240 112.980 41.695 ;
        RECT 106.195 40.995 112.980 41.240 ;
        RECT 110.840 39.360 111.440 39.610 ;
        RECT 101.650 39.220 111.440 39.360 ;
        RECT 110.840 38.970 111.440 39.220 ;
        RECT 83.430 37.125 83.590 37.265 ;
        RECT 56.175 36.265 69.740 36.965 ;
        RECT 56.175 35.985 56.875 36.265 ;
        RECT 55.860 35.855 56.875 35.985 ;
        RECT 44.900 35.245 45.800 35.575 ;
        RECT 44.400 34.945 45.800 35.245 ;
        RECT 54.155 35.155 56.875 35.855 ;
        RECT 55.860 35.025 56.760 35.155 ;
        RECT 44.400 31.200 44.700 34.945 ;
        RECT 44.900 34.615 45.800 34.945 ;
        RECT 57.080 34.365 58.210 35.535 ;
        RECT 69.040 34.070 69.740 36.265 ;
        RECT 72.495 36.145 73.075 36.340 ;
        RECT 83.430 36.145 83.570 37.125 ;
        RECT 72.495 36.005 83.570 36.145 ;
        RECT 70.920 34.725 72.050 35.895 ;
        RECT 72.495 35.700 73.075 36.005 ;
        RECT 68.940 33.110 69.840 34.070 ;
        RECT 46.225 31.895 47.355 33.065 ;
        RECT 47.590 31.200 48.490 31.890 ;
        RECT 57.080 31.320 58.210 32.490 ;
        RECT 44.400 31.060 48.490 31.200 ;
        RECT 44.400 28.960 44.700 31.060 ;
        RECT 47.590 30.930 48.490 31.060 ;
        RECT 44.900 28.960 45.800 29.290 ;
        RECT 44.400 28.660 45.800 28.960 ;
        RECT 44.400 25.090 44.700 28.660 ;
        RECT 44.900 28.330 45.800 28.660 ;
        RECT 46.260 25.800 47.390 26.970 ;
        RECT 47.590 25.090 48.490 25.485 ;
        RECT 44.400 24.790 48.490 25.090 ;
        RECT 41.845 24.525 42.745 24.745 ;
        RECT 45.200 23.215 45.500 24.790 ;
        RECT 47.590 24.525 48.490 24.790 ;
        RECT 44.900 22.255 45.800 23.215 ;
        RECT 36.090 19.375 37.220 20.545 ;
        RECT 46.215 19.395 47.345 20.565 ;
        RECT 95.300 17.525 96.430 18.695 ;
        RECT 138.180 14.655 140.550 16.985 ;
        RECT 138.580 8.815 140.150 10.345 ;
        RECT 128.250 6.605 129.820 8.135 ;
        RECT 106.315 4.685 107.885 6.215 ;
        RECT 83.975 3.020 85.545 4.550 ;
        RECT 61.800 1.480 63.370 3.010 ;
      LAYER met3 ;
        RECT 97.750 213.655 98.050 213.660 ;
        RECT 97.535 212.885 98.265 213.655 ;
        RECT 105.730 213.025 106.460 213.795 ;
        RECT 97.750 209.485 98.050 212.885 ;
        RECT 105.945 209.485 106.245 213.025 ;
        RECT 97.750 209.185 106.245 209.485 ;
        RECT 97.750 206.480 98.050 209.185 ;
        RECT 105.945 206.715 106.245 209.185 ;
        RECT 97.535 205.710 98.265 206.480 ;
        RECT 105.730 205.945 106.460 206.715 ;
        RECT 97.750 199.530 98.050 205.710 ;
        RECT 105.945 199.845 106.245 205.945 ;
        RECT 97.535 198.760 98.265 199.530 ;
        RECT 105.730 199.075 106.460 199.845 ;
        RECT 97.750 192.505 98.050 198.760 ;
        RECT 105.945 192.505 106.245 199.075 ;
        RECT 95.765 192.220 96.495 192.455 ;
        RECT 97.535 192.220 98.265 192.505 ;
        RECT 95.765 191.920 98.265 192.220 ;
        RECT 95.765 191.685 96.495 191.920 ;
        RECT 97.535 191.735 98.265 191.920 ;
        RECT 105.730 191.735 106.460 192.505 ;
        RECT 53.180 190.075 54.310 190.575 ;
        RECT 53.180 189.775 57.455 190.075 ;
        RECT 53.180 189.405 54.310 189.775 ;
        RECT 57.155 188.275 57.455 189.775 ;
        RECT 97.535 188.705 98.265 189.475 ;
        RECT 97.750 188.275 98.050 188.705 ;
        RECT 57.155 187.975 98.050 188.275 ;
        RECT 105.945 173.440 106.245 191.735 ;
        RECT 105.700 172.670 106.430 173.440 ;
        RECT 105.945 166.650 106.245 172.670 ;
        RECT 105.700 165.880 106.430 166.650 ;
        RECT 17.620 148.635 20.000 148.795 ;
        RECT 21.330 148.635 23.700 148.800 ;
        RECT 17.620 146.635 23.700 148.635 ;
        RECT 17.620 146.475 20.000 146.635 ;
        RECT 21.330 146.470 23.700 146.635 ;
        RECT 138.180 147.650 140.550 147.815 ;
        RECT 143.710 147.650 146.090 147.810 ;
        RECT 138.180 145.650 146.090 147.650 ;
        RECT 138.180 145.485 140.550 145.650 ;
        RECT 143.710 145.490 146.090 145.650 ;
        RECT 71.600 108.710 72.330 108.830 ;
        RECT 42.240 108.695 72.330 108.710 ;
        RECT 40.890 108.410 72.330 108.695 ;
        RECT 40.890 108.395 42.540 108.410 ;
        RECT 40.890 101.490 41.190 108.395 ;
        RECT 71.600 108.060 72.330 108.410 ;
        RECT 43.910 101.490 45.040 102.240 ;
        RECT 40.890 101.190 45.040 101.490 ;
        RECT 40.890 91.620 41.190 101.190 ;
        RECT 43.910 101.070 45.040 101.190 ;
        RECT 52.895 101.105 54.025 102.275 ;
        RECT 53.310 99.600 53.610 101.105 ;
        RECT 63.390 101.045 64.520 102.215 ;
        RECT 63.575 100.025 63.875 101.045 ;
        RECT 51.645 99.300 53.610 99.600 ;
        RECT 62.010 99.725 63.955 100.025 ;
        RECT 43.910 91.620 45.040 92.330 ;
        RECT 40.890 91.320 45.040 91.620 ;
        RECT 43.910 91.160 45.040 91.320 ;
        RECT 51.645 92.040 51.945 99.300 ;
        RECT 52.895 92.040 54.025 92.365 ;
        RECT 51.645 91.740 54.025 92.040 ;
        RECT 43.910 81.525 45.040 82.175 ;
        RECT 42.945 81.225 45.040 81.525 ;
        RECT 42.945 72.615 43.245 81.225 ;
        RECT 43.910 81.005 45.040 81.225 ;
        RECT 51.645 81.915 51.945 91.740 ;
        RECT 52.895 91.195 54.025 91.740 ;
        RECT 62.010 91.760 62.310 99.725 ;
        RECT 120.135 97.875 120.865 97.910 ;
        RECT 102.885 97.175 120.865 97.875 ;
        RECT 94.580 95.345 95.710 95.540 ;
        RECT 92.890 94.645 95.710 95.345 ;
        RECT 92.890 93.815 93.590 94.645 ;
        RECT 94.580 94.370 95.710 94.645 ;
        RECT 92.675 93.590 93.805 93.815 ;
        RECT 91.555 92.890 93.805 93.590 ;
        RECT 102.885 93.130 103.585 97.175 ;
        RECT 120.135 97.140 120.865 97.175 ;
        RECT 112.910 95.345 114.040 95.540 ;
        RECT 111.220 94.645 114.040 95.345 ;
        RECT 111.220 93.815 111.920 94.645 ;
        RECT 112.910 94.370 114.040 94.645 ;
        RECT 111.005 93.590 112.135 93.815 ;
        RECT 63.390 91.760 64.520 92.320 ;
        RECT 91.555 92.250 92.255 92.890 ;
        RECT 92.675 92.645 93.805 92.890 ;
        RECT 91.555 92.235 92.775 92.250 ;
        RECT 62.010 91.460 64.520 91.760 ;
        RECT 52.895 81.915 54.025 82.350 ;
        RECT 51.645 81.615 54.025 81.915 ;
        RECT 50.465 75.770 51.195 76.005 ;
        RECT 51.645 75.770 51.945 81.615 ;
        RECT 52.895 81.180 54.025 81.615 ;
        RECT 62.010 82.010 62.310 91.460 ;
        RECT 63.390 91.150 64.520 91.460 ;
        RECT 89.510 91.535 92.775 92.235 ;
        RECT 102.710 91.960 103.840 93.130 ;
        RECT 109.970 92.890 112.135 93.590 ;
        RECT 109.970 92.320 110.670 92.890 ;
        RECT 111.005 92.645 112.135 92.890 ;
        RECT 107.840 92.250 110.890 92.320 ;
        RECT 89.510 90.745 90.210 91.535 ;
        RECT 91.645 91.080 92.775 91.535 ;
        RECT 107.840 91.620 111.105 92.250 ;
        RECT 107.840 90.745 108.540 91.620 ;
        RECT 109.975 91.080 111.105 91.620 ;
        RECT 89.295 90.365 90.425 90.745 ;
        RECT 107.625 90.450 108.755 90.745 ;
        RECT 86.340 89.665 90.425 90.365 ;
        RECT 86.340 88.585 87.040 89.665 ;
        RECT 89.295 89.575 90.425 89.665 ;
        RECT 104.670 89.750 108.755 90.450 ;
        RECT 104.670 88.605 105.370 89.750 ;
        RECT 107.625 89.575 108.755 89.750 ;
        RECT 86.080 87.415 87.210 88.585 ;
        RECT 104.410 87.435 105.540 88.605 ;
        RECT 86.355 85.830 87.055 87.415 ;
        RECT 88.615 85.830 89.745 86.205 ;
        RECT 86.355 85.130 89.745 85.830 ;
        RECT 104.685 85.970 105.385 87.435 ;
        RECT 106.945 85.970 108.075 86.205 ;
        RECT 104.685 85.270 108.075 85.970 ;
        RECT 88.615 85.035 89.745 85.130 ;
        RECT 106.945 85.035 108.075 85.270 ;
        RECT 88.970 84.055 89.670 85.035 ;
        RECT 90.690 84.055 91.820 84.780 ;
        RECT 88.970 83.610 91.820 84.055 ;
        RECT 107.300 84.195 108.000 85.035 ;
        RECT 109.020 84.195 110.150 84.780 ;
        RECT 107.300 83.610 110.150 84.195 ;
        RECT 88.970 83.355 91.605 83.610 ;
        RECT 107.300 83.495 109.935 83.610 ;
        RECT 90.905 82.835 91.605 83.355 ;
        RECT 109.235 82.835 109.935 83.495 ;
        RECT 63.390 82.010 64.520 82.465 ;
        RECT 72.435 82.215 73.565 82.615 ;
        RECT 62.010 81.710 64.520 82.010 ;
        RECT 50.465 75.470 51.945 75.770 ;
        RECT 50.465 75.235 51.195 75.470 ;
        RECT 43.910 72.735 45.040 73.170 ;
        RECT 51.645 73.035 51.945 75.470 ;
        RECT 52.895 73.045 54.025 73.145 ;
        RECT 62.010 73.045 62.310 81.710 ;
        RECT 63.390 81.295 64.520 81.710 ;
        RECT 70.885 81.915 73.565 82.215 ;
        RECT 63.390 73.045 64.520 73.290 ;
        RECT 52.895 73.035 64.520 73.045 ;
        RECT 51.645 72.745 64.520 73.035 ;
        RECT 51.645 72.735 54.025 72.745 ;
        RECT 43.910 72.615 51.945 72.735 ;
        RECT 42.945 72.435 51.945 72.615 ;
        RECT 42.945 72.315 45.040 72.435 ;
        RECT 43.910 72.000 45.040 72.315 ;
        RECT 52.895 71.975 54.025 72.735 ;
        RECT 63.390 72.120 64.520 72.745 ;
        RECT 70.885 72.525 71.185 81.915 ;
        RECT 72.435 81.445 73.565 81.915 ;
        RECT 90.690 81.665 91.820 82.835 ;
        RECT 109.020 81.665 110.150 82.835 ;
        RECT 90.770 80.920 91.470 81.665 ;
        RECT 92.960 80.920 94.090 81.295 ;
        RECT 90.770 80.220 94.090 80.920 ;
        RECT 92.960 80.125 94.090 80.220 ;
        RECT 96.115 80.940 97.245 81.295 ;
        RECT 109.100 80.940 109.800 81.665 ;
        RECT 111.290 80.940 112.420 81.295 ;
        RECT 96.115 80.240 112.420 80.940 ;
        RECT 96.115 80.125 97.245 80.240 ;
        RECT 93.175 79.800 93.875 80.125 ;
        RECT 96.340 79.800 97.040 80.125 ;
        RECT 93.175 79.100 97.040 79.800 ;
        RECT 94.340 77.055 95.470 77.250 ;
        RECT 92.600 76.355 95.470 77.055 ;
        RECT 92.600 75.525 93.300 76.355 ;
        RECT 94.340 76.080 95.470 76.355 ;
        RECT 92.385 75.300 93.515 75.525 ;
        RECT 91.370 74.600 93.515 75.300 ;
        RECT 91.370 74.090 92.070 74.600 ;
        RECT 92.385 74.355 93.515 74.600 ;
        RECT 89.025 73.960 92.075 74.090 ;
        RECT 89.025 73.390 92.485 73.960 ;
        RECT 72.030 72.525 73.160 72.990 ;
        RECT 70.885 72.225 73.160 72.525 ;
        RECT 89.025 72.455 89.725 73.390 ;
        RECT 91.355 72.790 92.485 73.390 ;
        RECT 70.885 71.675 71.185 72.225 ;
        RECT 72.030 71.820 73.160 72.225 ;
        RECT 89.005 72.220 90.135 72.455 ;
        RECT 48.615 71.375 71.185 71.675 ;
        RECT 85.855 71.520 90.135 72.220 ;
        RECT 48.615 65.535 48.915 71.375 ;
        RECT 56.570 69.110 56.870 71.375 ;
        RECT 85.855 70.315 86.555 71.520 ;
        RECT 89.005 71.285 90.135 71.520 ;
        RECT 85.790 69.145 86.920 70.315 ;
        RECT 56.385 68.340 57.115 69.110 ;
        RECT 85.855 67.450 86.555 69.145 ;
        RECT 88.325 67.450 89.455 67.915 ;
        RECT 85.855 66.750 89.455 67.450 ;
        RECT 88.325 66.745 89.455 66.750 ;
        RECT 49.505 65.535 50.635 65.970 ;
        RECT 48.615 65.235 50.635 65.535 ;
        RECT 45.945 58.795 46.675 59.075 ;
        RECT 48.615 58.795 48.915 65.235 ;
        RECT 49.505 64.800 50.635 65.235 ;
        RECT 88.680 65.675 89.380 66.745 ;
        RECT 90.400 65.675 91.530 66.490 ;
        RECT 88.680 65.320 91.530 65.675 ;
        RECT 88.680 64.975 91.315 65.320 ;
        RECT 90.615 64.545 91.315 64.975 ;
        RECT 90.400 63.375 91.530 64.545 ;
        RECT 90.480 62.540 91.180 63.375 ;
        RECT 92.670 62.540 93.800 63.005 ;
        RECT 90.480 61.840 93.800 62.540 ;
        RECT 92.670 61.835 93.800 61.840 ;
        RECT 95.825 62.305 96.955 63.005 ;
        RECT 101.445 62.305 102.145 80.240 ;
        RECT 111.290 80.125 112.420 80.240 ;
        RECT 114.445 80.125 115.575 81.295 ;
        RECT 111.635 79.820 112.335 80.125 ;
        RECT 114.660 79.820 115.360 80.125 ;
        RECT 111.635 79.120 115.360 79.820 ;
        RECT 112.940 76.810 114.070 77.005 ;
        RECT 111.250 76.110 114.070 76.810 ;
        RECT 111.250 75.280 111.950 76.110 ;
        RECT 112.940 75.835 114.070 76.110 ;
        RECT 111.035 75.055 112.165 75.280 ;
        RECT 109.995 74.355 112.165 75.055 ;
        RECT 109.995 73.845 110.695 74.355 ;
        RECT 111.035 74.110 112.165 74.355 ;
        RECT 107.655 73.715 110.705 73.845 ;
        RECT 107.655 73.145 111.135 73.715 ;
        RECT 107.655 72.210 108.355 73.145 ;
        RECT 109.995 73.130 111.135 73.145 ;
        RECT 110.005 72.545 111.135 73.130 ;
        RECT 107.655 71.975 108.785 72.210 ;
        RECT 104.485 71.275 108.785 71.975 ;
        RECT 104.485 70.085 105.185 71.275 ;
        RECT 107.655 71.040 108.785 71.275 ;
        RECT 104.440 68.915 105.570 70.085 ;
        RECT 104.485 67.435 105.185 68.915 ;
        RECT 106.975 67.435 108.105 67.670 ;
        RECT 104.485 66.735 108.105 67.435 ;
        RECT 106.975 66.500 108.105 66.735 ;
        RECT 107.330 65.660 108.030 66.500 ;
        RECT 109.050 65.660 110.180 66.245 ;
        RECT 107.330 65.075 110.180 65.660 ;
        RECT 107.330 64.960 109.965 65.075 ;
        RECT 109.265 64.300 109.965 64.960 ;
        RECT 109.050 63.130 110.180 64.300 ;
        RECT 109.130 62.305 109.830 63.130 ;
        RECT 111.320 62.305 112.450 62.760 ;
        RECT 95.825 61.835 112.450 62.305 ;
        RECT 92.885 61.420 93.585 61.835 ;
        RECT 96.040 61.605 112.450 61.835 ;
        RECT 96.040 61.420 96.750 61.605 ;
        RECT 92.885 60.720 96.750 61.420 ;
        RECT 100.555 60.940 101.255 61.605 ;
        RECT 111.320 61.590 112.450 61.605 ;
        RECT 114.475 61.590 115.605 62.760 ;
        RECT 111.535 61.185 112.235 61.590 ;
        RECT 114.700 61.185 115.400 61.590 ;
        RECT 100.555 60.200 101.330 60.940 ;
        RECT 111.535 60.485 115.400 61.185 ;
        RECT 100.610 60.160 101.330 60.200 ;
        RECT 49.505 58.795 50.635 59.280 ;
        RECT 45.945 58.495 50.635 58.795 ;
        RECT 45.945 58.305 46.675 58.495 ;
        RECT 49.505 58.110 50.635 58.495 ;
        RECT 103.320 58.910 107.990 58.940 ;
        RECT 103.320 58.240 110.590 58.910 ;
        RECT 103.320 55.495 104.020 58.240 ;
        RECT 106.910 58.210 110.590 58.240 ;
        RECT 106.910 57.125 107.610 58.210 ;
        RECT 109.890 57.125 110.590 58.210 ;
        RECT 106.675 55.955 107.805 57.125 ;
        RECT 109.675 55.955 110.805 57.125 ;
        RECT 104.425 55.495 105.555 55.715 ;
        RECT 70.960 54.150 72.080 55.330 ;
        RECT 102.125 54.795 105.555 55.495 ;
        RECT 102.125 53.605 102.825 54.795 ;
        RECT 104.425 54.545 105.555 54.795 ;
        RECT 104.090 53.605 105.220 54.040 ;
        RECT 102.125 53.305 105.220 53.605 ;
        RECT 49.505 52.180 50.635 52.615 ;
        RECT 48.605 51.880 50.635 52.180 ;
        RECT 48.605 45.700 48.905 51.880 ;
        RECT 49.505 51.445 50.635 51.880 ;
        RECT 59.520 49.555 60.650 50.725 ;
        RECT 70.960 50.400 72.080 51.580 ;
        RECT 102.125 50.565 102.825 53.305 ;
        RECT 104.090 52.870 105.220 53.305 ;
        RECT 102.125 49.985 102.890 50.565 ;
        RECT 104.090 49.985 105.220 50.420 ;
        RECT 102.125 49.865 105.220 49.985 ;
        RECT 58.005 48.230 59.135 49.400 ;
        RECT 59.935 48.840 60.235 49.555 ;
        RECT 58.545 46.685 58.845 48.230 ;
        RECT 59.520 47.670 60.650 48.840 ;
        RECT 71.055 48.670 72.185 49.840 ;
        RECT 102.185 49.685 105.220 49.865 ;
        RECT 59.935 47.015 60.235 47.670 ;
        RECT 71.520 47.270 71.820 48.670 ;
        RECT 59.520 46.685 60.650 47.015 ;
        RECT 58.545 46.385 60.650 46.685 ;
        RECT 49.505 45.790 50.635 45.990 ;
        RECT 58.545 45.790 58.845 46.385 ;
        RECT 59.520 45.845 60.650 46.385 ;
        RECT 70.995 46.100 72.125 47.270 ;
        RECT 49.505 45.700 58.845 45.790 ;
        RECT 48.605 45.490 58.845 45.700 ;
        RECT 48.605 45.400 50.635 45.490 ;
        RECT 49.505 44.820 50.635 45.400 ;
        RECT 59.935 45.140 60.235 45.845 ;
        RECT 59.520 43.970 60.650 45.140 ;
        RECT 71.520 44.765 71.820 46.100 ;
        RECT 102.185 44.830 102.885 49.685 ;
        RECT 104.090 49.250 105.220 49.685 ;
        RECT 104.090 46.435 105.220 46.670 ;
        RECT 103.745 45.500 105.220 46.435 ;
        RECT 103.745 44.830 104.445 45.500 ;
        RECT 104.765 44.830 105.895 45.065 ;
        RECT 59.935 43.320 60.235 43.970 ;
        RECT 71.105 43.595 72.235 44.765 ;
        RECT 102.185 44.130 105.895 44.830 ;
        RECT 59.520 42.150 60.650 43.320 ;
        RECT 71.520 42.155 71.820 43.595 ;
        RECT 59.935 41.580 60.235 42.150 ;
        RECT 59.520 40.410 60.650 41.580 ;
        RECT 71.105 40.985 72.235 42.155 ;
        RECT 103.745 41.745 104.445 44.130 ;
        RECT 104.765 43.895 105.895 44.130 ;
        RECT 107.175 42.405 108.305 43.575 ;
        RECT 109.905 42.445 111.035 43.615 ;
        RECT 103.745 41.445 104.585 41.745 ;
        RECT 35.040 39.325 36.680 39.355 ;
        RECT 37.430 39.325 38.560 39.760 ;
        RECT 46.240 39.335 47.370 39.770 ;
        RECT 59.935 39.745 60.235 40.410 ;
        RECT 35.040 39.025 38.560 39.325 ;
        RECT 35.040 32.855 35.340 39.025 ;
        RECT 37.430 38.590 38.560 39.025 ;
        RECT 44.065 39.035 47.370 39.335 ;
        RECT 37.080 32.855 38.210 33.055 ;
        RECT 35.040 32.555 38.210 32.855 ;
        RECT 17.620 29.555 20.000 29.715 ;
        RECT 21.330 29.555 23.700 29.720 ;
        RECT 17.620 27.555 23.700 29.555 ;
        RECT 17.620 27.395 20.000 27.555 ;
        RECT 21.330 27.390 23.700 27.555 ;
        RECT 35.040 26.635 35.340 32.555 ;
        RECT 37.080 31.885 38.210 32.555 ;
        RECT 44.065 32.640 44.365 39.035 ;
        RECT 46.240 38.600 47.370 39.035 ;
        RECT 59.520 38.575 60.650 39.745 ;
        RECT 71.520 39.670 71.820 40.985 ;
        RECT 104.085 40.855 104.385 41.445 ;
        RECT 107.390 40.855 108.090 42.405 ;
        RECT 110.105 40.855 110.805 42.445 ;
        RECT 95.410 40.155 110.805 40.855 ;
        RECT 71.105 38.500 72.235 39.670 ;
        RECT 71.520 37.785 71.820 38.500 ;
        RECT 71.190 37.015 71.920 37.785 ;
        RECT 57.080 35.100 58.210 35.535 ;
        RECT 70.920 35.100 72.050 35.895 ;
        RECT 54.265 34.800 72.050 35.100 ;
        RECT 46.225 32.695 47.355 33.065 ;
        RECT 54.265 32.695 54.565 34.800 ;
        RECT 57.080 34.365 58.210 34.800 ;
        RECT 70.920 34.725 72.050 34.800 ;
        RECT 44.065 32.630 45.250 32.640 ;
        RECT 46.225 32.630 54.565 32.695 ;
        RECT 44.065 32.395 54.565 32.630 ;
        RECT 44.065 32.330 47.355 32.395 ;
        RECT 37.080 26.635 38.210 26.940 ;
        RECT 35.040 26.335 38.210 26.635 ;
        RECT 35.040 20.110 35.340 26.335 ;
        RECT 37.080 25.770 38.210 26.335 ;
        RECT 44.065 26.605 44.365 32.330 ;
        RECT 46.225 31.895 47.355 32.330 ;
        RECT 55.895 32.055 56.615 32.180 ;
        RECT 57.080 32.055 58.210 32.490 ;
        RECT 55.895 31.755 58.210 32.055 ;
        RECT 55.895 31.400 56.615 31.755 ;
        RECT 57.080 31.320 58.210 31.755 ;
        RECT 46.260 26.605 47.390 26.970 ;
        RECT 44.065 26.305 47.390 26.605 ;
        RECT 36.090 20.110 37.220 20.545 ;
        RECT 35.040 20.025 37.220 20.110 ;
        RECT 44.065 20.025 44.365 26.305 ;
        RECT 44.995 26.285 45.295 26.305 ;
        RECT 46.260 25.800 47.390 26.305 ;
        RECT 46.215 20.025 47.345 20.565 ;
        RECT 35.040 19.810 47.345 20.025 ;
        RECT 36.090 19.725 47.345 19.810 ;
        RECT 36.090 19.375 37.220 19.725 ;
        RECT 46.215 19.395 47.345 19.725 ;
        RECT 95.410 18.695 96.110 40.155 ;
        RECT 95.300 18.460 96.430 18.695 ;
        RECT 100.100 18.460 122.555 34.760 ;
        RECT 95.300 17.760 122.555 18.460 ;
        RECT 95.300 17.525 96.430 17.760 ;
        RECT 100.100 12.310 122.555 17.760 ;
        RECT 138.180 16.820 140.550 16.985 ;
        RECT 143.710 16.820 146.090 16.980 ;
        RECT 138.180 14.820 146.090 16.820 ;
        RECT 138.180 14.655 140.550 14.820 ;
        RECT 143.710 14.660 146.090 14.820 ;
        RECT 139.365 10.345 144.940 10.580 ;
        RECT 138.580 10.340 144.940 10.345 ;
        RECT 138.580 8.820 145.690 10.340 ;
        RECT 138.580 8.815 144.940 8.820 ;
        RECT 139.365 8.580 144.940 8.815 ;
        RECT 128.250 8.130 134.610 8.370 ;
        RECT 128.250 6.610 135.360 8.130 ;
        RECT 106.315 6.210 112.675 6.450 ;
        RECT 128.250 6.370 134.610 6.610 ;
        RECT 83.975 4.545 90.335 4.785 ;
        RECT 106.315 4.690 113.425 6.210 ;
        RECT 67.330 3.020 68.910 3.040 ;
        RECT 61.800 2.020 68.910 3.020 ;
        RECT 83.975 3.025 91.085 4.545 ;
        RECT 106.315 4.450 112.675 4.690 ;
        RECT 83.975 2.785 90.335 3.025 ;
        RECT 61.800 1.480 63.370 2.020 ;
        RECT 67.330 1.520 68.910 2.020 ;
      LAYER met4 ;
        RECT 3.490 224.760 3.990 225.055 ;
        RECT 4.290 224.760 7.670 225.055 ;
        RECT 7.970 224.760 11.350 225.055 ;
        RECT 11.650 224.760 15.030 225.055 ;
        RECT 15.330 224.760 18.710 225.055 ;
        RECT 19.010 224.760 22.390 225.055 ;
        RECT 22.690 224.760 26.070 225.055 ;
        RECT 26.370 224.760 29.750 225.055 ;
        RECT 30.050 224.760 33.430 225.055 ;
        RECT 33.730 224.760 37.110 225.055 ;
        RECT 37.410 224.760 40.790 225.055 ;
        RECT 41.090 224.760 44.470 225.055 ;
        RECT 44.770 224.760 48.150 225.055 ;
        RECT 48.450 224.760 51.830 225.055 ;
        RECT 52.130 224.760 55.510 225.055 ;
        RECT 55.810 224.760 59.190 225.055 ;
        RECT 59.490 224.760 62.870 225.055 ;
        RECT 63.170 224.760 66.550 225.055 ;
        RECT 66.850 224.760 70.230 225.055 ;
        RECT 70.530 224.760 73.910 225.055 ;
        RECT 74.210 224.760 77.590 225.055 ;
        RECT 77.890 224.760 81.270 225.055 ;
        RECT 81.570 224.760 84.950 225.055 ;
        RECT 85.250 224.760 88.630 225.055 ;
        RECT 3.490 224.755 88.770 224.760 ;
        RECT 3.490 148.655 5.490 224.755 ;
        RECT 17.645 148.655 19.975 148.800 ;
        RECT 3.490 146.655 20.085 148.655 ;
        RECT 143.735 147.670 146.065 147.815 ;
        RECT 158.355 147.670 160.355 224.150 ;
        RECT 3.490 29.575 5.490 146.655 ;
        RECT 17.645 146.470 19.975 146.655 ;
        RECT 143.735 145.670 160.355 147.670 ;
        RECT 143.735 145.485 146.065 145.670 ;
        RECT 100.605 60.185 101.335 60.915 ;
        RECT 56.070 54.285 57.700 55.510 ;
        RECT 56.070 54.275 57.065 54.285 ;
        RECT 57.075 54.275 57.700 54.285 ;
        RECT 56.070 53.050 57.700 54.275 ;
        RECT 70.955 54.175 72.085 55.305 ;
        RECT 71.370 52.270 71.670 54.175 ;
        RECT 57.570 51.970 71.670 52.270 ;
        RECT 57.570 43.745 57.870 51.970 ;
        RECT 71.370 51.555 71.670 51.970 ;
        RECT 70.955 50.425 72.085 51.555 ;
        RECT 55.950 43.725 57.870 43.745 ;
        RECT 54.935 43.445 57.870 43.725 ;
        RECT 54.935 43.425 56.250 43.445 ;
        RECT 54.935 31.940 55.235 43.425 ;
        RECT 100.620 34.620 101.320 60.185 ;
        RECT 55.890 31.940 56.620 32.155 ;
        RECT 54.935 31.640 56.620 31.940 ;
        RECT 55.890 31.425 56.620 31.640 ;
        RECT 17.645 29.575 19.975 29.720 ;
        RECT 3.490 27.575 20.085 29.575 ;
        RECT 3.490 1.005 5.490 27.575 ;
        RECT 17.645 27.390 19.975 27.575 ;
        RECT 100.240 12.450 122.415 34.620 ;
        RECT 143.735 16.840 146.065 16.985 ;
        RECT 158.355 16.840 160.355 145.670 ;
        RECT 143.735 14.840 160.355 16.840 ;
        RECT 143.735 14.655 146.065 14.840 ;
        RECT 144.900 10.345 157.735 10.580 ;
        RECT 144.135 8.815 157.735 10.345 ;
        RECT 144.900 8.580 157.735 8.815 ;
        RECT 133.805 6.605 135.335 8.135 ;
        RECT 111.870 4.685 113.400 6.215 ;
        RECT 89.530 4.280 91.060 4.550 ;
        RECT 67.355 2.950 68.885 3.045 ;
        RECT 89.530 3.020 91.160 4.280 ;
        RECT 67.355 1.515 69.015 2.950 ;
        RECT 68.015 1.000 69.015 1.515 ;
        RECT 68.015 0.670 68.240 1.000 ;
        RECT 68.840 0.670 69.015 1.000 ;
        RECT 90.160 1.000 91.160 3.020 ;
        RECT 90.160 0.830 90.320 1.000 ;
        RECT 90.920 0.830 91.160 1.000 ;
        RECT 112.140 1.000 113.140 4.685 ;
        RECT 112.140 0.495 112.400 1.000 ;
        RECT 113.000 0.495 113.140 1.000 ;
        RECT 134.290 1.000 135.290 6.605 ;
        RECT 134.290 0.790 134.480 1.000 ;
        RECT 135.080 0.790 135.290 1.000 ;
        RECT 155.735 1.000 157.735 8.580 ;
        RECT 158.355 1.005 160.355 14.840 ;
        RECT 155.735 0.670 156.560 1.000 ;
        RECT 157.160 0.670 157.735 1.000 ;
  END
END tt_um_Burrows_Katie
END LIBRARY

