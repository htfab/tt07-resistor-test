VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Burrows_Katie
  CLASS BLOCK ;
  FOREIGN tt_um_Burrow_Katie ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNADIFFAREA 17.639999 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 4.410000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 4.410000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 6.095000 ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNAGATEAREA 4.000000 ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 158.360 0.260 160.360 224.145 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3.490 0.200 5.490 225.040 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 52.415 209.310 53.085 209.390 ;
        RECT 52.415 206.520 58.355 209.310 ;
      LAYER nwell ;
        RECT 97.890 207.500 104.310 212.780 ;
        RECT 105.970 207.500 112.390 212.780 ;
      LAYER pwell ;
        RECT 52.415 206.440 53.085 206.520 ;
        RECT 52.415 204.610 53.085 204.690 ;
        RECT 52.415 201.820 58.355 204.610 ;
      LAYER nwell ;
        RECT 63.075 203.430 65.495 206.710 ;
        RECT 92.055 203.465 94.475 206.745 ;
      LAYER pwell ;
        RECT 52.415 201.740 53.085 201.820 ;
      LAYER nwell ;
        RECT 97.890 200.510 104.310 205.790 ;
        RECT 105.970 200.510 112.390 205.790 ;
      LAYER pwell ;
        RECT 52.415 198.075 53.085 198.155 ;
        RECT 52.415 195.285 58.355 198.075 ;
        RECT 52.415 195.205 53.085 195.285 ;
      LAYER nwell ;
        RECT 76.600 194.120 83.020 199.400 ;
        RECT 97.890 193.520 104.310 198.800 ;
        RECT 105.970 193.520 112.390 198.800 ;
      LAYER pwell ;
        RECT 52.415 193.265 53.085 193.345 ;
        RECT 52.415 190.475 58.355 193.265 ;
        RECT 52.415 190.395 53.085 190.475 ;
      LAYER nwell ;
        RECT 76.600 187.205 83.020 192.485 ;
        RECT 97.890 186.495 104.310 191.775 ;
        RECT 105.970 186.495 112.390 191.775 ;
      LAYER pwell ;
        RECT 45.320 184.870 45.990 184.950 ;
        RECT 45.320 182.080 53.260 184.870 ;
        RECT 45.320 182.000 45.990 182.080 ;
        RECT 45.320 180.395 45.990 180.475 ;
        RECT 45.320 177.605 53.260 180.395 ;
        RECT 45.320 177.525 45.990 177.605 ;
        RECT 45.320 175.780 45.990 175.860 ;
        RECT 45.320 172.990 53.260 175.780 ;
        RECT 45.320 172.910 45.990 172.990 ;
        RECT 45.300 170.205 45.970 170.285 ;
        RECT 45.300 167.415 53.240 170.205 ;
      LAYER nwell ;
        RECT 88.450 169.495 90.870 172.775 ;
        RECT 106.195 167.880 112.615 173.160 ;
      LAYER pwell ;
        RECT 45.300 167.335 45.970 167.415 ;
        RECT 45.300 165.690 45.970 165.770 ;
        RECT 45.300 162.900 53.240 165.690 ;
        RECT 45.300 162.820 45.970 162.900 ;
        RECT 45.300 161.100 45.970 161.180 ;
        RECT 45.300 158.310 53.240 161.100 ;
      LAYER nwell ;
        RECT 88.445 159.495 90.865 162.775 ;
        RECT 106.195 160.770 112.615 166.050 ;
      LAYER pwell ;
        RECT 45.300 158.230 45.970 158.310 ;
        RECT 45.250 108.400 45.920 108.480 ;
        RECT 45.250 103.610 51.190 108.400 ;
        RECT 45.250 103.530 45.920 103.610 ;
      LAYER nwell ;
        RECT 54.515 103.420 60.935 108.700 ;
        RECT 64.665 103.420 71.085 108.700 ;
        RECT 73.945 103.375 80.365 108.655 ;
      LAYER pwell ;
        RECT 45.250 98.585 45.920 98.665 ;
        RECT 45.250 93.795 51.190 98.585 ;
        RECT 45.250 93.715 45.920 93.795 ;
      LAYER nwell ;
        RECT 54.515 93.525 60.935 98.805 ;
        RECT 64.665 93.545 71.085 98.825 ;
        RECT 73.945 93.485 80.365 98.765 ;
      LAYER pwell ;
        RECT 45.250 88.425 45.920 88.505 ;
        RECT 45.250 83.635 51.190 88.425 ;
        RECT 45.250 83.555 45.920 83.635 ;
      LAYER nwell ;
        RECT 54.515 83.480 60.935 88.760 ;
        RECT 64.665 83.605 71.085 88.885 ;
        RECT 73.900 83.650 80.320 88.930 ;
        RECT 97.345 82.390 103.765 95.360 ;
        RECT 115.690 82.390 122.110 95.360 ;
      LAYER pwell ;
        RECT 45.250 79.360 45.920 79.440 ;
        RECT 45.250 74.570 51.190 79.360 ;
        RECT 45.250 74.490 45.920 74.570 ;
      LAYER nwell ;
        RECT 54.515 74.280 60.935 79.560 ;
        RECT 64.665 74.185 71.085 79.465 ;
        RECT 73.945 74.090 80.365 79.370 ;
      LAYER pwell ;
        RECT 50.935 71.145 51.605 71.225 ;
        RECT 50.935 67.355 57.875 71.145 ;
        RECT 50.935 67.275 51.605 67.355 ;
        RECT 50.935 64.455 51.605 64.535 ;
        RECT 50.935 60.665 57.875 64.455 ;
        RECT 50.935 60.585 51.605 60.665 ;
        RECT 50.935 57.765 51.605 57.845 ;
        RECT 50.935 53.975 57.875 57.765 ;
      LAYER nwell ;
        RECT 63.860 55.625 72.280 69.365 ;
        RECT 76.215 56.045 84.635 69.845 ;
        RECT 97.040 64.100 103.460 77.070 ;
        RECT 115.695 63.855 122.115 76.825 ;
      LAYER pwell ;
        RECT 50.935 53.895 51.605 53.975 ;
        RECT 50.935 51.125 51.605 51.205 ;
        RECT 50.935 47.335 57.875 51.125 ;
        RECT 50.935 47.255 51.605 47.335 ;
        RECT 37.465 44.925 38.135 45.005 ;
        RECT 47.590 44.925 48.260 45.005 ;
        RECT 37.465 41.135 44.505 44.925 ;
        RECT 47.590 41.135 54.630 44.925 ;
        RECT 37.465 41.055 38.135 41.135 ;
        RECT 47.590 41.055 48.260 41.135 ;
      LAYER nwell ;
        RECT 64.115 38.920 72.535 52.660 ;
        RECT 76.235 38.400 84.655 52.200 ;
        RECT 112.880 44.825 121.300 57.165 ;
      LAYER pwell ;
        RECT 37.465 38.230 38.135 38.310 ;
        RECT 47.590 38.230 48.260 38.310 ;
        RECT 37.465 34.440 44.505 38.230 ;
        RECT 47.590 34.440 54.630 38.230 ;
        RECT 71.945 35.470 72.615 35.550 ;
        RECT 58.495 35.295 59.165 35.375 ;
        RECT 37.465 34.360 38.135 34.440 ;
        RECT 47.590 34.360 48.260 34.440 ;
        RECT 58.495 33.875 66.435 35.295 ;
        RECT 71.945 34.050 79.885 35.470 ;
        RECT 71.945 33.970 72.615 34.050 ;
        RECT 58.495 33.795 59.165 33.875 ;
        RECT 37.465 32.115 38.135 32.195 ;
        RECT 47.590 32.115 48.260 32.195 ;
        RECT 37.465 28.325 44.505 32.115 ;
        RECT 47.590 28.325 54.630 32.115 ;
        RECT 37.465 28.245 38.135 28.325 ;
        RECT 47.590 28.245 48.260 28.325 ;
        RECT 37.465 25.710 38.135 25.790 ;
        RECT 47.590 25.710 48.260 25.790 ;
        RECT 37.465 21.920 44.505 25.710 ;
        RECT 47.590 21.920 54.630 25.710 ;
        RECT 37.465 21.840 38.135 21.920 ;
        RECT 47.590 21.840 48.260 21.920 ;
      LAYER li1 ;
        RECT 98.765 212.760 99.295 213.290 ;
        RECT 107.045 212.760 107.575 213.290 ;
        RECT 98.880 212.365 99.180 212.760 ;
        RECT 98.575 212.195 103.325 212.365 ;
        RECT 103.760 211.700 104.090 212.445 ;
        RECT 107.160 212.365 107.460 212.760 ;
        RECT 106.655 212.195 111.405 212.365 ;
        RECT 104.375 211.700 104.905 211.835 ;
        RECT 103.760 211.370 104.905 211.700 ;
        RECT 52.585 208.395 52.915 209.220 ;
        RECT 53.620 209.140 54.320 210.330 ;
        RECT 97.370 210.100 97.970 210.700 ;
        RECT 53.350 208.970 58.100 209.140 ;
        RECT 51.675 207.695 52.915 208.395 ;
        RECT 52.585 206.610 52.915 207.695 ;
        RECT 58.780 207.550 59.310 208.080 ;
        RECT 98.575 207.915 103.325 208.085 ;
        RECT 103.010 207.500 103.180 207.915 ;
        RECT 103.760 207.835 104.090 211.370 ;
        RECT 104.375 211.305 104.905 211.370 ;
        RECT 111.840 211.545 112.170 212.445 ;
        RECT 112.475 211.545 113.005 211.685 ;
        RECT 111.840 211.215 113.005 211.545 ;
        RECT 105.565 210.240 106.165 210.840 ;
        RECT 106.655 207.915 111.405 208.085 ;
        RECT 106.860 207.770 107.165 207.915 ;
        RECT 111.840 207.835 112.170 211.215 ;
        RECT 112.475 211.155 113.005 211.215 ;
        RECT 106.865 207.500 107.165 207.770 ;
        RECT 53.350 206.690 58.100 206.860 ;
        RECT 63.880 206.760 64.410 207.290 ;
        RECT 92.965 206.760 93.495 207.290 ;
        RECT 102.830 206.970 103.360 207.500 ;
        RECT 106.750 206.970 107.280 207.500 ;
        RECT 53.420 206.360 53.720 206.690 ;
        RECT 53.305 205.830 53.835 206.360 ;
        RECT 63.995 206.295 64.165 206.760 ;
        RECT 64.965 206.375 65.295 206.395 ;
        RECT 63.800 206.125 64.470 206.295 ;
        RECT 52.585 203.495 52.915 204.520 ;
        RECT 53.610 204.440 54.310 205.265 ;
        RECT 62.340 205.050 63.230 205.940 ;
        RECT 53.350 204.270 58.100 204.440 ;
        RECT 63.800 203.950 64.470 204.015 ;
        RECT 51.675 202.795 52.915 203.495 ;
        RECT 63.785 203.845 64.470 203.950 ;
        RECT 63.785 203.485 64.185 203.845 ;
        RECT 64.945 203.765 65.295 206.375 ;
        RECT 93.090 206.330 93.390 206.760 ;
        RECT 92.780 206.160 93.450 206.330 ;
        RECT 93.090 206.125 93.390 206.160 ;
        RECT 91.250 205.050 92.140 205.940 ;
        RECT 92.780 203.880 93.450 204.050 ;
        RECT 93.925 203.940 94.255 206.410 ;
        RECT 98.765 205.565 99.295 206.095 ;
        RECT 107.045 205.565 107.575 206.095 ;
        RECT 98.880 205.375 99.180 205.565 ;
        RECT 98.575 205.205 103.325 205.375 ;
        RECT 58.780 202.895 59.310 203.425 ;
        RECT 63.700 202.955 64.230 203.485 ;
        RECT 52.585 201.910 52.915 202.795 ;
        RECT 64.965 202.410 65.295 203.765 ;
        RECT 93.090 203.505 93.390 203.880 ;
        RECT 93.900 203.800 94.255 203.940 ;
        RECT 103.760 204.780 104.090 205.455 ;
        RECT 107.160 205.375 107.460 205.565 ;
        RECT 106.655 205.205 111.405 205.375 ;
        RECT 104.395 204.780 104.925 204.920 ;
        RECT 103.760 204.450 104.925 204.780 ;
        RECT 92.965 202.975 93.495 203.505 ;
        RECT 93.900 202.505 94.230 203.800 ;
        RECT 97.370 202.925 97.970 203.525 ;
        RECT 53.350 201.990 58.100 202.160 ;
        RECT 53.380 201.550 53.680 201.990 ;
        RECT 64.965 201.980 65.505 202.410 ;
        RECT 64.975 201.880 65.505 201.980 ;
        RECT 93.775 201.975 94.305 202.505 ;
        RECT 53.265 201.020 53.795 201.550 ;
        RECT 98.575 200.925 103.325 201.095 ;
        RECT 103.095 200.435 103.265 200.925 ;
        RECT 103.760 200.845 104.090 204.450 ;
        RECT 104.395 204.390 104.925 204.450 ;
        RECT 111.840 204.780 112.170 205.455 ;
        RECT 112.475 204.780 113.005 204.920 ;
        RECT 111.840 204.450 113.005 204.780 ;
        RECT 105.565 203.160 106.165 203.760 ;
        RECT 106.655 200.925 111.405 201.095 ;
        RECT 106.950 200.435 107.250 200.925 ;
        RECT 111.840 200.845 112.170 204.450 ;
        RECT 112.475 204.390 113.005 204.450 ;
        RECT 81.245 198.985 81.945 200.205 ;
        RECT 102.915 199.905 103.445 200.435 ;
        RECT 106.835 199.905 107.365 200.435 ;
        RECT 52.585 196.960 52.915 197.985 ;
        RECT 53.535 197.905 54.235 198.835 ;
        RECT 77.285 198.815 82.035 198.985 ;
        RECT 82.470 198.945 82.800 199.065 ;
        RECT 82.470 198.245 83.770 198.945 ;
        RECT 98.765 198.590 99.295 199.120 ;
        RECT 107.045 198.660 107.575 199.190 ;
        RECT 98.880 198.385 99.180 198.590 ;
        RECT 53.350 197.735 58.100 197.905 ;
        RECT 51.675 196.260 52.915 196.960 ;
        RECT 58.780 196.500 59.310 197.030 ;
        RECT 76.045 196.515 76.575 197.045 ;
        RECT 52.585 195.375 52.915 196.260 ;
        RECT 53.350 195.455 58.100 195.625 ;
        RECT 53.435 195.130 53.735 195.455 ;
        RECT 53.320 194.600 53.850 195.130 ;
        RECT 77.285 194.535 82.035 194.705 ;
        RECT 77.605 194.150 77.905 194.535 ;
        RECT 82.470 194.455 82.800 198.245 ;
        RECT 98.575 198.215 103.325 198.385 ;
        RECT 103.760 197.605 104.090 198.465 ;
        RECT 107.160 198.385 107.460 198.660 ;
        RECT 106.655 198.215 111.405 198.385 ;
        RECT 104.395 197.605 104.925 197.810 ;
        RECT 103.760 197.280 104.925 197.605 ;
        RECT 111.840 197.605 112.170 198.465 ;
        RECT 112.475 197.605 113.005 197.810 ;
        RECT 111.840 197.280 113.005 197.605 ;
        RECT 103.760 197.275 104.825 197.280 ;
        RECT 111.840 197.275 112.905 197.280 ;
        RECT 97.370 195.975 97.970 196.575 ;
        RECT 52.585 192.270 52.915 193.175 ;
        RECT 53.590 193.095 54.290 193.910 ;
        RECT 77.490 193.620 78.020 194.150 ;
        RECT 98.575 193.935 103.325 194.105 ;
        RECT 103.095 193.555 103.265 193.935 ;
        RECT 103.760 193.855 104.090 197.275 ;
        RECT 105.565 196.290 106.165 196.890 ;
        RECT 106.655 193.935 111.405 194.105 ;
        RECT 106.950 193.555 107.250 193.935 ;
        RECT 111.840 193.855 112.170 197.275 ;
        RECT 53.350 192.925 58.100 193.095 ;
        RECT 51.675 191.570 52.915 192.270 ;
        RECT 81.245 192.070 81.945 193.100 ;
        RECT 102.915 193.025 103.445 193.555 ;
        RECT 106.835 193.025 107.365 193.555 ;
        RECT 52.585 190.565 52.915 191.570 ;
        RECT 58.780 191.455 59.310 191.985 ;
        RECT 77.285 191.900 82.035 192.070 ;
        RECT 82.470 192.050 82.800 192.150 ;
        RECT 82.470 191.350 83.770 192.050 ;
        RECT 98.765 191.615 99.295 192.145 ;
        RECT 107.045 191.680 107.575 192.210 ;
        RECT 98.945 191.360 99.115 191.615 ;
        RECT 53.350 190.645 58.100 190.815 ;
        RECT 53.400 190.310 53.700 190.645 ;
        RECT 53.320 189.780 53.850 190.310 ;
        RECT 76.025 189.240 76.555 189.770 ;
        RECT 77.285 187.620 82.035 187.790 ;
        RECT 77.605 187.285 77.905 187.620 ;
        RECT 82.470 187.540 82.800 191.350 ;
        RECT 98.575 191.190 103.325 191.360 ;
        RECT 103.760 190.505 104.090 191.440 ;
        RECT 107.160 191.360 107.460 191.680 ;
        RECT 106.655 191.190 111.405 191.360 ;
        RECT 104.395 190.505 104.925 190.745 ;
        RECT 103.760 190.215 104.925 190.505 ;
        RECT 103.760 190.175 104.825 190.215 ;
        RECT 97.370 188.950 97.970 189.550 ;
        RECT 77.490 186.755 78.020 187.285 ;
        RECT 98.575 186.910 103.325 187.080 ;
        RECT 103.095 186.395 103.265 186.910 ;
        RECT 103.760 186.830 104.090 190.175 ;
        RECT 111.840 190.065 112.170 191.440 ;
        RECT 112.475 190.065 113.005 190.305 ;
        RECT 111.840 189.775 113.005 190.065 ;
        RECT 111.840 189.735 112.905 189.775 ;
        RECT 105.565 188.950 106.165 189.550 ;
        RECT 106.655 186.910 111.405 187.080 ;
        RECT 106.950 186.395 107.250 186.910 ;
        RECT 111.840 186.830 112.170 189.735 ;
        RECT 45.490 184.700 45.820 184.780 ;
        RECT 46.355 184.700 47.055 185.875 ;
        RECT 102.915 185.865 103.445 186.395 ;
        RECT 106.835 185.865 107.365 186.395 ;
        RECT 44.430 184.000 45.820 184.700 ;
        RECT 46.235 184.530 53.025 184.700 ;
        RECT 45.490 182.170 45.820 184.000 ;
        RECT 53.640 183.185 54.170 183.715 ;
        RECT 46.235 182.250 53.025 182.420 ;
        RECT 52.720 181.890 53.020 182.250 ;
        RECT 52.630 181.360 53.160 181.890 ;
        RECT 58.325 181.170 58.495 183.050 ;
        RECT 118.660 182.380 118.830 183.050 ;
        RECT 45.490 180.245 45.820 180.305 ;
        RECT 44.430 179.545 45.820 180.245 ;
        RECT 46.355 180.225 47.055 181.145 ;
        RECT 46.235 180.055 53.025 180.225 ;
        RECT 45.490 177.695 45.820 179.545 ;
        RECT 53.640 178.730 54.170 179.260 ;
        RECT 58.325 178.750 58.495 180.630 ;
        RECT 118.660 179.960 118.830 181.840 ;
        RECT 46.235 177.775 53.025 177.945 ;
        RECT 52.715 177.375 53.015 177.775 ;
        RECT 52.630 176.845 53.160 177.375 ;
        RECT 45.490 175.645 45.820 175.690 ;
        RECT 44.430 174.945 45.820 175.645 ;
        RECT 46.355 175.610 47.055 176.580 ;
        RECT 58.325 176.330 58.495 178.210 ;
        RECT 118.660 177.540 118.830 179.420 ;
        RECT 118.660 176.330 118.830 177.000 ;
        RECT 46.235 175.440 53.025 175.610 ;
        RECT 45.490 173.080 45.820 174.945 ;
        RECT 53.640 174.035 54.170 174.565 ;
        RECT 46.235 173.160 53.025 173.330 ;
        RECT 52.720 172.775 53.020 173.160 ;
        RECT 52.630 172.245 53.160 172.775 ;
        RECT 89.030 172.745 89.560 173.275 ;
        RECT 106.780 172.745 107.480 173.765 ;
        RECT 89.175 172.360 89.475 172.745 ;
        RECT 106.780 172.640 111.630 172.745 ;
        RECT 106.880 172.575 111.630 172.640 ;
        RECT 89.175 172.190 89.845 172.360 ;
        RECT 89.175 172.130 89.475 172.190 ;
        RECT 45.470 170.100 45.800 170.115 ;
        RECT 44.430 169.400 45.800 170.100 ;
        RECT 46.270 170.035 46.970 171.010 ;
        RECT 87.675 170.740 88.565 171.630 ;
        RECT 90.320 171.385 90.650 172.440 ;
        RECT 112.065 172.085 112.395 172.825 ;
        RECT 112.065 171.385 113.510 172.085 ;
        RECT 90.320 170.685 91.585 171.385 ;
        RECT 46.215 169.865 53.005 170.035 ;
        RECT 89.175 169.910 89.845 170.080 ;
        RECT 45.470 167.505 45.800 169.400 ;
        RECT 89.175 169.305 89.475 169.910 ;
        RECT 90.320 169.830 90.650 170.685 ;
        RECT 105.535 169.885 106.135 170.485 ;
        RECT 53.615 168.325 54.145 168.855 ;
        RECT 89.055 168.775 89.585 169.305 ;
        RECT 106.980 168.465 107.680 168.475 ;
        RECT 106.880 168.295 111.630 168.465 ;
        RECT 46.215 167.585 53.005 167.755 ;
        RECT 45.470 165.460 45.800 165.600 ;
        RECT 46.270 165.520 46.970 166.560 ;
        RECT 52.285 166.550 52.985 167.585 ;
        RECT 106.980 167.350 107.680 168.295 ;
        RECT 112.065 168.215 112.395 171.385 ;
        RECT 106.780 165.635 107.480 166.595 ;
        RECT 106.780 165.545 111.630 165.635 ;
        RECT 44.495 164.760 45.800 165.460 ;
        RECT 46.215 165.350 53.005 165.520 ;
        RECT 106.880 165.465 111.630 165.545 ;
        RECT 112.065 165.530 112.395 165.715 ;
        RECT 45.470 162.990 45.800 164.760 ;
        RECT 112.065 164.830 113.420 165.530 ;
        RECT 53.645 164.015 54.175 164.545 ;
        RECT 46.215 163.070 53.005 163.240 ;
        RECT 52.285 162.010 52.985 163.070 ;
        RECT 89.045 162.685 89.575 163.215 ;
        RECT 93.770 162.715 94.300 163.245 ;
        RECT 105.535 163.095 106.135 163.695 ;
        RECT 89.180 162.360 89.480 162.685 ;
        RECT 89.170 162.190 89.840 162.360 ;
        RECT 89.180 162.120 89.480 162.190 ;
        RECT 45.470 160.995 45.800 161.010 ;
        RECT 44.430 160.295 45.800 160.995 ;
        RECT 46.270 160.930 46.970 161.985 ;
        RECT 46.215 160.760 53.005 160.930 ;
        RECT 87.765 160.780 88.655 161.670 ;
        RECT 90.315 161.430 90.645 162.440 ;
        RECT 45.470 158.400 45.800 160.295 ;
        RECT 90.315 160.730 91.650 161.430 ;
        RECT 106.880 161.185 111.630 161.355 ;
        RECT 53.625 159.415 54.155 159.945 ;
        RECT 89.170 159.910 89.840 160.080 ;
        RECT 89.180 159.315 89.480 159.910 ;
        RECT 90.315 159.830 90.645 160.730 ;
        RECT 106.980 160.210 107.680 161.185 ;
        RECT 112.065 161.105 112.395 164.830 ;
        RECT 89.055 158.785 89.585 159.315 ;
        RECT 46.215 158.480 53.005 158.650 ;
        RECT 52.265 157.260 52.965 158.480 ;
        RECT 45.685 153.510 45.855 155.390 ;
        RECT 110.690 154.720 110.860 155.390 ;
        RECT 45.685 151.090 45.855 152.970 ;
        RECT 110.690 152.300 110.860 154.180 ;
        RECT 45.685 148.670 45.855 150.550 ;
        RECT 110.690 149.880 110.860 151.760 ;
        RECT 45.685 146.250 45.855 148.130 ;
        RECT 110.690 147.460 110.860 149.340 ;
        RECT 45.685 143.830 45.855 145.710 ;
        RECT 110.690 145.040 110.860 146.920 ;
        RECT 45.685 141.410 45.855 143.290 ;
        RECT 110.690 142.620 110.860 144.500 ;
        RECT 45.685 138.990 45.855 140.870 ;
        RECT 110.690 140.200 110.860 142.080 ;
        RECT 45.685 136.570 45.855 138.450 ;
        RECT 110.690 137.780 110.860 139.660 ;
        RECT 110.690 136.570 110.860 137.240 ;
        RECT 46.055 108.910 46.585 109.080 ;
        RECT 55.040 108.920 55.570 109.090 ;
        RECT 65.275 108.920 65.805 109.090 ;
        RECT 45.420 107.065 45.750 108.310 ;
        RECT 46.230 108.230 46.400 108.910 ;
        RECT 55.215 108.285 55.385 108.920 ;
        RECT 46.185 108.060 50.935 108.230 ;
        RECT 55.200 108.115 59.950 108.285 ;
        RECT 46.230 108.055 46.400 108.060 ;
        RECT 44.065 106.065 45.750 107.065 ;
        RECT 60.385 106.490 60.715 108.365 ;
        RECT 65.450 108.285 65.620 108.920 ;
        RECT 65.350 108.115 70.100 108.285 ;
        RECT 70.535 106.530 70.865 108.365 ;
        RECT 78.665 108.240 79.365 109.670 ;
        RECT 74.630 108.070 79.380 108.240 ;
        RECT 78.665 108.060 79.365 108.070 ;
        RECT 45.420 103.700 45.750 106.065 ;
        RECT 51.595 105.925 52.125 106.455 ;
        RECT 60.385 106.420 61.760 106.490 ;
        RECT 70.535 106.420 71.970 106.530 ;
        RECT 60.385 106.250 62.045 106.420 ;
        RECT 70.535 106.250 72.070 106.420 ;
        RECT 60.385 106.160 61.760 106.250 ;
        RECT 70.535 106.200 71.970 106.250 ;
        RECT 54.035 103.960 54.565 104.490 ;
        RECT 46.185 103.780 50.935 103.950 ;
        RECT 55.200 103.835 59.950 104.005 ;
        RECT 46.255 103.330 46.425 103.780 ;
        RECT 55.240 103.365 55.410 103.835 ;
        RECT 60.385 103.755 60.715 106.160 ;
        RECT 64.195 103.930 64.725 104.460 ;
        RECT 65.350 103.835 70.100 104.005 ;
        RECT 45.795 102.330 46.795 103.330 ;
        RECT 54.780 102.365 55.780 103.365 ;
        RECT 65.735 103.305 65.905 103.835 ;
        RECT 70.535 103.755 70.865 106.200 ;
        RECT 73.395 105.720 73.925 106.250 ;
        RECT 74.630 103.790 79.380 103.960 ;
        RECT 65.275 102.305 66.275 103.305 ;
        RECT 74.650 103.285 74.820 103.790 ;
        RECT 74.245 102.395 75.135 103.285 ;
        RECT 79.815 102.750 80.145 108.320 ;
        RECT 82.970 104.425 83.140 105.095 ;
        RECT 79.530 102.705 80.145 102.750 ;
        RECT 79.430 102.535 80.145 102.705 ;
        RECT 79.530 102.420 80.145 102.535 ;
        RECT 82.970 102.005 83.140 103.885 ;
        RECT 123.805 103.215 123.975 105.095 ;
        RECT 46.055 100.060 46.585 100.230 ;
        RECT 45.420 97.270 45.750 98.495 ;
        RECT 46.230 98.415 46.400 100.060 ;
        RECT 55.040 98.960 55.570 99.130 ;
        RECT 65.275 98.980 65.805 99.150 ;
        RECT 46.185 98.245 50.935 98.415 ;
        RECT 55.215 98.390 55.385 98.960 ;
        RECT 55.200 98.220 59.950 98.390 ;
        RECT 44.065 96.270 45.750 97.270 ;
        RECT 45.420 93.885 45.750 96.270 ;
        RECT 51.615 95.815 52.145 96.345 ;
        RECT 60.385 96.100 60.715 98.470 ;
        RECT 65.450 98.410 65.620 98.980 ;
        RECT 64.195 97.735 64.725 98.265 ;
        RECT 65.350 98.240 70.100 98.410 ;
        RECT 70.535 96.205 70.865 98.490 ;
        RECT 78.665 98.350 79.365 99.765 ;
        RECT 82.970 99.585 83.140 101.465 ;
        RECT 123.805 100.795 123.975 102.675 ;
        RECT 123.805 99.585 123.975 100.255 ;
        RECT 74.630 98.180 79.380 98.350 ;
        RECT 78.665 98.155 79.365 98.180 ;
        RECT 60.385 96.070 61.805 96.100 ;
        RECT 70.535 96.070 71.970 96.205 ;
        RECT 60.385 95.900 62.045 96.070 ;
        RECT 70.535 95.900 72.070 96.070 ;
        RECT 60.385 95.770 61.805 95.900 ;
        RECT 70.535 95.875 71.970 95.900 ;
        RECT 46.185 93.965 50.935 94.135 ;
        RECT 54.035 94.030 54.565 94.560 ;
        RECT 46.255 93.420 46.425 93.965 ;
        RECT 55.200 93.940 59.950 94.110 ;
        RECT 55.240 93.455 55.410 93.940 ;
        RECT 60.385 93.860 60.715 95.770 ;
        RECT 65.350 93.960 70.100 94.130 ;
        RECT 45.795 92.420 46.795 93.420 ;
        RECT 54.780 92.455 55.780 93.455 ;
        RECT 65.735 93.410 65.905 93.960 ;
        RECT 70.535 93.880 70.865 95.875 ;
        RECT 73.415 95.755 73.945 96.285 ;
        RECT 74.630 93.900 79.380 94.070 ;
        RECT 65.275 92.410 66.275 93.410 ;
        RECT 74.650 93.385 74.820 93.900 ;
        RECT 74.245 92.495 75.135 93.385 ;
        RECT 79.815 93.235 80.145 98.430 ;
        RECT 93.260 95.695 93.790 96.225 ;
        RECT 96.465 95.630 97.465 96.630 ;
        RECT 112.295 96.290 112.825 96.820 ;
        RECT 98.155 95.850 98.685 96.020 ;
        RECT 94.560 93.930 95.560 94.905 ;
        RECT 96.225 94.745 96.755 94.770 ;
        RECT 96.225 94.600 96.840 94.745 ;
        RECT 96.595 94.575 96.840 94.600 ;
        RECT 94.560 93.905 96.400 93.930 ;
        RECT 95.135 93.760 96.400 93.905 ;
        RECT 79.530 93.185 80.145 93.235 ;
        RECT 79.430 93.015 80.145 93.185 ;
        RECT 79.530 92.905 80.145 93.015 ;
        RECT 93.530 92.340 94.530 93.340 ;
        RECT 96.230 93.270 96.400 93.760 ;
        RECT 96.670 93.685 96.840 94.575 ;
        RECT 97.190 94.305 97.360 95.630 ;
        RECT 98.335 94.945 98.505 95.850 ;
        RECT 114.795 95.630 115.795 96.630 ;
        RECT 116.485 95.850 117.015 96.020 ;
        RECT 98.030 94.775 102.780 94.945 ;
        RECT 98.030 94.305 102.780 94.315 ;
        RECT 97.190 94.145 102.780 94.305 ;
        RECT 97.190 94.135 98.160 94.145 ;
        RECT 103.215 93.780 103.545 95.025 ;
        RECT 104.595 93.780 105.595 94.220 ;
        RECT 112.890 93.930 113.890 94.905 ;
        RECT 114.555 94.745 115.085 94.770 ;
        RECT 114.555 94.600 115.170 94.745 ;
        RECT 114.925 94.575 115.170 94.600 ;
        RECT 112.890 93.905 114.730 93.930 ;
        RECT 96.670 93.515 102.780 93.685 ;
        RECT 103.215 93.450 105.595 93.780 ;
        RECT 113.465 93.760 114.730 93.905 ;
        RECT 96.230 93.100 97.730 93.270 ;
        RECT 95.175 92.930 95.790 93.100 ;
        RECT 95.620 92.865 95.790 92.930 ;
        RECT 97.560 93.055 97.730 93.100 ;
        RECT 97.560 92.885 102.780 93.055 ;
        RECT 95.620 92.695 97.270 92.865 ;
        RECT 97.100 92.625 97.270 92.695 ;
        RECT 97.100 92.455 97.745 92.625 ;
        RECT 94.360 92.235 94.530 92.340 ;
        RECT 97.575 92.425 97.745 92.455 ;
        RECT 97.575 92.255 102.780 92.425 ;
        RECT 94.360 92.065 97.165 92.235 ;
        RECT 91.180 90.835 92.180 91.835 ;
        RECT 96.995 91.795 97.165 92.065 ;
        RECT 93.420 91.585 96.805 91.755 ;
        RECT 96.995 91.625 102.780 91.795 ;
        RECT 93.420 91.520 93.590 91.585 ;
        RECT 93.060 91.350 93.590 91.520 ;
        RECT 94.215 91.060 96.080 91.230 ;
        RECT 89.860 90.620 90.390 90.705 ;
        RECT 89.860 90.450 90.650 90.620 ;
        RECT 90.480 90.050 90.650 90.450 ;
        RECT 91.830 90.510 92.000 90.835 ;
        RECT 94.215 90.510 94.385 91.060 ;
        RECT 91.830 90.340 94.385 90.510 ;
        RECT 95.910 90.535 96.080 91.060 ;
        RECT 96.635 91.165 96.805 91.585 ;
        RECT 96.635 90.995 102.780 91.165 ;
        RECT 95.910 90.365 102.780 90.535 ;
        RECT 91.470 90.050 93.745 90.075 ;
        RECT 55.040 89.190 55.570 89.360 ;
        RECT 65.275 89.315 65.805 89.485 ;
        RECT 46.055 88.840 46.585 89.010 ;
        RECT 45.420 87.910 45.750 88.335 ;
        RECT 46.230 88.255 46.400 88.840 ;
        RECT 55.225 88.345 55.395 89.190 ;
        RECT 65.460 88.470 65.630 89.315 ;
        RECT 46.185 88.085 50.935 88.255 ;
        RECT 55.200 88.175 59.950 88.345 ;
        RECT 44.065 86.910 45.750 87.910 ;
        RECT 45.420 83.725 45.750 86.910 ;
        RECT 51.595 85.740 52.125 86.270 ;
        RECT 60.385 86.115 60.715 88.425 ;
        RECT 65.350 88.300 70.100 88.470 ;
        RECT 64.195 87.730 64.725 88.260 ;
        RECT 70.535 86.265 70.865 88.550 ;
        RECT 78.615 88.515 79.315 89.955 ;
        RECT 90.480 89.905 93.745 90.050 ;
        RECT 90.480 89.880 91.640 89.905 ;
        RECT 93.575 89.735 102.780 89.905 ;
        RECT 87.965 89.275 88.965 89.675 ;
        RECT 87.965 89.105 102.780 89.275 ;
        RECT 87.965 88.675 88.965 89.105 ;
        RECT 98.030 88.615 102.780 88.645 ;
        RECT 74.585 88.345 79.335 88.515 ;
        RECT 70.535 86.210 71.970 86.265 ;
        RECT 60.385 86.050 61.850 86.115 ;
        RECT 60.385 85.880 62.045 86.050 ;
        RECT 70.535 86.040 72.070 86.210 ;
        RECT 70.535 85.935 71.970 86.040 ;
        RECT 73.355 85.995 73.885 86.525 ;
        RECT 60.385 85.785 61.850 85.880 ;
        RECT 54.035 83.980 54.565 84.510 ;
        RECT 46.185 83.805 50.935 83.975 ;
        RECT 55.200 83.895 59.950 84.065 ;
        RECT 46.255 83.265 46.425 83.805 ;
        RECT 55.240 83.440 55.410 83.895 ;
        RECT 60.385 83.815 60.715 85.785 ;
        RECT 65.350 84.020 70.100 84.190 ;
        RECT 65.735 83.555 65.905 84.020 ;
        RECT 70.535 83.940 70.865 85.935 ;
        RECT 74.585 84.065 79.335 84.235 ;
        RECT 74.590 83.705 74.760 84.065 ;
        RECT 45.795 82.265 46.795 83.265 ;
        RECT 54.780 82.440 55.780 83.440 ;
        RECT 65.275 82.555 66.275 83.555 ;
        RECT 74.320 82.705 75.320 83.705 ;
        RECT 79.770 82.830 80.100 88.595 ;
        RECT 96.490 88.475 102.780 88.615 ;
        RECT 96.490 88.445 98.245 88.475 ;
        RECT 96.490 88.345 96.660 88.445 ;
        RECT 89.860 88.175 96.660 88.345 ;
        RECT 97.055 88.015 98.195 88.030 ;
        RECT 97.055 87.860 102.780 88.015 ;
        RECT 97.055 87.810 97.225 87.860 ;
        RECT 98.030 87.845 102.780 87.860 ;
        RECT 90.915 87.640 97.225 87.810 ;
        RECT 90.915 87.295 91.085 87.640 ;
        RECT 98.030 87.365 102.780 87.385 ;
        RECT 97.515 87.325 102.780 87.365 ;
        RECT 90.500 86.295 91.500 87.295 ;
        RECT 92.640 87.215 102.780 87.325 ;
        RECT 92.640 87.195 98.185 87.215 ;
        RECT 92.640 87.155 97.685 87.195 ;
        RECT 92.640 86.880 92.810 87.155 ;
        RECT 92.195 86.710 92.810 86.880 ;
        RECT 93.295 86.585 102.780 86.755 ;
        RECT 93.295 85.870 93.465 86.585 ;
        RECT 94.760 85.955 102.780 86.125 ;
        RECT 92.575 84.870 93.575 85.870 ;
        RECT 94.760 85.360 94.930 85.955 ;
        RECT 94.300 85.190 94.930 85.360 ;
        RECT 94.480 85.150 94.930 85.190 ;
        RECT 95.470 85.325 102.780 85.495 ;
        RECT 95.470 84.455 95.640 85.325 ;
        RECT 93.450 84.285 95.640 84.455 ;
        RECT 96.080 84.695 102.780 84.865 ;
        RECT 93.450 83.925 93.620 84.285 ;
        RECT 92.575 83.340 93.620 83.925 ;
        RECT 96.080 83.605 96.250 84.695 ;
        RECT 94.685 83.535 96.250 83.605 ;
        RECT 94.505 83.435 96.250 83.535 ;
        RECT 96.700 84.065 102.780 84.235 ;
        RECT 94.505 83.365 95.035 83.435 ;
        RECT 92.575 82.925 93.575 83.340 ;
        RECT 96.700 83.050 96.870 84.065 ;
        RECT 79.395 82.665 80.100 82.830 ;
        RECT 95.640 82.880 96.870 83.050 ;
        RECT 97.190 83.435 102.780 83.605 ;
        RECT 79.395 82.660 79.925 82.665 ;
        RECT 95.640 82.385 95.810 82.880 ;
        RECT 94.845 81.385 95.845 82.385 ;
        RECT 97.190 82.110 97.360 83.435 ;
        RECT 98.030 82.805 102.780 82.975 ;
        RECT 98.415 82.385 98.585 82.805 ;
        RECT 103.215 82.725 103.545 93.450 ;
        RECT 104.595 93.220 105.595 93.450 ;
        RECT 111.860 92.340 112.860 93.340 ;
        RECT 114.560 93.270 114.730 93.760 ;
        RECT 115.000 93.685 115.170 94.575 ;
        RECT 115.520 94.305 115.690 95.630 ;
        RECT 116.665 94.945 116.835 95.850 ;
        RECT 116.375 94.775 121.125 94.945 ;
        RECT 116.375 94.305 121.125 94.315 ;
        RECT 115.520 94.145 121.125 94.305 ;
        RECT 115.520 94.135 116.490 94.145 ;
        RECT 115.000 93.515 121.125 93.685 ;
        RECT 114.560 93.100 116.060 93.270 ;
        RECT 113.505 92.930 114.120 93.100 ;
        RECT 113.950 92.865 114.120 92.930 ;
        RECT 115.890 93.055 116.060 93.100 ;
        RECT 115.890 92.885 121.125 93.055 ;
        RECT 113.950 92.695 115.600 92.865 ;
        RECT 115.430 92.625 115.600 92.695 ;
        RECT 115.430 92.455 116.075 92.625 ;
        RECT 112.690 92.235 112.860 92.340 ;
        RECT 115.905 92.425 116.075 92.455 ;
        RECT 115.905 92.255 121.125 92.425 ;
        RECT 112.690 92.065 115.495 92.235 ;
        RECT 109.510 90.835 110.510 91.835 ;
        RECT 115.325 91.795 115.495 92.065 ;
        RECT 111.750 91.585 115.135 91.755 ;
        RECT 115.325 91.625 121.125 91.795 ;
        RECT 111.750 91.520 111.920 91.585 ;
        RECT 111.390 91.350 111.920 91.520 ;
        RECT 112.545 91.060 114.410 91.230 ;
        RECT 108.190 90.620 108.720 90.705 ;
        RECT 108.190 90.450 108.980 90.620 ;
        RECT 108.810 90.050 108.980 90.450 ;
        RECT 110.160 90.510 110.330 90.835 ;
        RECT 112.545 90.510 112.715 91.060 ;
        RECT 110.160 90.340 112.715 90.510 ;
        RECT 114.240 90.535 114.410 91.060 ;
        RECT 114.965 91.165 115.135 91.585 ;
        RECT 114.965 90.995 121.125 91.165 ;
        RECT 114.240 90.365 121.125 90.535 ;
        RECT 109.800 90.050 112.075 90.075 ;
        RECT 108.810 89.905 112.075 90.050 ;
        RECT 108.810 89.880 109.970 89.905 ;
        RECT 111.905 89.735 121.125 89.905 ;
        RECT 106.295 89.275 107.295 89.695 ;
        RECT 121.560 89.650 121.890 95.025 ;
        RECT 106.295 89.105 121.125 89.275 ;
        RECT 106.295 88.695 107.295 89.105 ;
        RECT 121.560 88.950 123.005 89.650 ;
        RECT 116.375 88.615 121.125 88.645 ;
        RECT 114.820 88.475 121.125 88.615 ;
        RECT 114.820 88.445 116.575 88.475 ;
        RECT 114.820 88.345 114.990 88.445 ;
        RECT 108.190 88.175 114.990 88.345 ;
        RECT 115.385 88.015 116.525 88.030 ;
        RECT 115.385 87.860 121.125 88.015 ;
        RECT 115.385 87.810 115.555 87.860 ;
        RECT 116.375 87.845 121.125 87.860 ;
        RECT 109.245 87.640 115.555 87.810 ;
        RECT 109.245 87.295 109.415 87.640 ;
        RECT 116.375 87.365 121.125 87.385 ;
        RECT 115.845 87.325 121.125 87.365 ;
        RECT 108.830 86.295 109.830 87.295 ;
        RECT 110.970 87.215 121.125 87.325 ;
        RECT 110.970 87.195 116.515 87.215 ;
        RECT 110.970 87.155 116.015 87.195 ;
        RECT 110.970 86.880 111.140 87.155 ;
        RECT 110.525 86.710 111.140 86.880 ;
        RECT 111.625 86.585 121.125 86.755 ;
        RECT 111.625 85.870 111.795 86.585 ;
        RECT 113.090 85.955 121.125 86.125 ;
        RECT 110.905 84.870 111.905 85.870 ;
        RECT 113.090 85.360 113.260 85.955 ;
        RECT 112.630 85.190 113.260 85.360 ;
        RECT 112.810 85.150 113.260 85.190 ;
        RECT 113.800 85.325 121.125 85.495 ;
        RECT 113.800 84.455 113.970 85.325 ;
        RECT 111.780 84.285 113.970 84.455 ;
        RECT 114.410 84.695 121.125 84.865 ;
        RECT 111.780 83.925 111.950 84.285 ;
        RECT 110.905 83.340 111.950 83.925 ;
        RECT 114.410 83.605 114.580 84.695 ;
        RECT 113.015 83.535 114.580 83.605 ;
        RECT 112.835 83.435 114.580 83.535 ;
        RECT 115.030 84.065 121.125 84.235 ;
        RECT 112.835 83.365 113.365 83.435 ;
        RECT 110.905 82.925 111.905 83.340 ;
        RECT 115.030 83.050 115.200 84.065 ;
        RECT 113.970 82.880 115.200 83.050 ;
        RECT 115.520 83.435 121.125 83.605 ;
        RECT 113.970 82.385 114.140 82.880 ;
        RECT 96.765 82.075 97.360 82.110 ;
        RECT 96.585 81.940 97.360 82.075 ;
        RECT 96.585 81.905 97.115 81.940 ;
        RECT 98.000 81.385 99.000 82.385 ;
        RECT 113.175 81.385 114.175 82.385 ;
        RECT 115.520 82.110 115.690 83.435 ;
        RECT 116.375 82.805 121.125 82.975 ;
        RECT 116.745 82.385 116.915 82.805 ;
        RECT 121.560 82.725 121.890 88.950 ;
        RECT 115.095 82.075 115.690 82.110 ;
        RECT 114.915 81.940 115.690 82.075 ;
        RECT 114.915 81.905 115.445 81.940 ;
        RECT 116.330 81.385 117.330 82.385 ;
        RECT 46.055 79.765 46.585 79.935 ;
        RECT 45.420 77.340 45.750 79.270 ;
        RECT 46.230 79.190 46.400 79.765 ;
        RECT 55.040 79.755 55.570 79.925 ;
        RECT 65.275 79.800 65.805 79.970 ;
        RECT 46.185 79.020 50.935 79.190 ;
        RECT 55.215 79.145 55.385 79.755 ;
        RECT 54.035 78.560 54.565 79.090 ;
        RECT 55.200 78.975 59.950 79.145 ;
        RECT 43.695 76.340 45.750 77.340 ;
        RECT 60.385 77.165 60.715 79.225 ;
        RECT 65.450 79.050 65.620 79.800 ;
        RECT 78.865 79.655 79.395 79.660 ;
        RECT 78.685 79.490 79.395 79.655 ;
        RECT 64.195 78.465 64.725 78.995 ;
        RECT 65.350 78.880 70.100 79.050 ;
        RECT 60.385 77.115 61.815 77.165 ;
        RECT 51.615 76.540 52.145 77.070 ;
        RECT 60.385 76.945 62.045 77.115 ;
        RECT 60.385 76.835 61.815 76.945 ;
        RECT 70.535 76.935 70.865 79.130 ;
        RECT 78.685 78.955 79.385 79.490 ;
        RECT 74.630 78.785 79.385 78.955 ;
        RECT 78.685 78.770 79.385 78.785 ;
        RECT 70.535 76.885 71.745 76.935 ;
        RECT 45.420 74.660 45.750 76.340 ;
        RECT 46.185 74.740 50.935 74.910 ;
        RECT 46.255 74.260 46.425 74.740 ;
        RECT 55.200 74.695 59.950 74.865 ;
        RECT 45.795 73.260 46.795 74.260 ;
        RECT 55.240 74.235 55.410 74.695 ;
        RECT 60.385 74.615 60.715 76.835 ;
        RECT 70.535 76.715 72.070 76.885 ;
        RECT 70.535 76.605 71.745 76.715 ;
        RECT 65.350 74.600 70.100 74.770 ;
        RECT 65.735 74.380 65.905 74.600 ;
        RECT 70.535 74.520 70.865 76.605 ;
        RECT 73.375 76.295 73.905 76.825 ;
        RECT 74.640 74.675 74.810 74.695 ;
        RECT 74.630 74.505 79.380 74.675 ;
        RECT 54.780 73.235 55.780 74.235 ;
        RECT 65.275 73.380 66.275 74.380 ;
        RECT 74.640 74.080 74.810 74.505 ;
        RECT 73.915 73.080 74.915 74.080 ;
        RECT 79.815 73.390 80.145 79.035 ;
        RECT 92.950 77.310 93.480 77.840 ;
        RECT 96.225 77.340 97.225 78.340 ;
        RECT 97.865 77.560 98.395 77.730 ;
        RECT 94.270 75.640 95.270 76.615 ;
        RECT 95.935 76.455 96.465 76.480 ;
        RECT 95.935 76.310 96.550 76.455 ;
        RECT 96.305 76.285 96.550 76.310 ;
        RECT 94.270 75.615 96.110 75.640 ;
        RECT 94.845 75.470 96.110 75.615 ;
        RECT 93.240 74.050 94.240 75.050 ;
        RECT 95.940 74.980 96.110 75.470 ;
        RECT 96.380 75.395 96.550 76.285 ;
        RECT 96.900 76.015 97.070 77.340 ;
        RECT 98.045 76.655 98.215 77.560 ;
        RECT 111.600 76.935 112.130 77.465 ;
        RECT 114.825 77.095 115.825 78.095 ;
        RECT 116.515 77.315 117.045 77.485 ;
        RECT 97.725 76.485 102.475 76.655 ;
        RECT 97.725 76.015 102.475 76.025 ;
        RECT 96.900 75.855 102.475 76.015 ;
        RECT 96.900 75.845 97.870 75.855 ;
        RECT 96.380 75.225 102.475 75.395 ;
        RECT 95.940 74.810 97.440 74.980 ;
        RECT 94.885 74.640 95.500 74.810 ;
        RECT 95.330 74.575 95.500 74.640 ;
        RECT 97.270 74.765 97.440 74.810 ;
        RECT 97.270 74.595 102.475 74.765 ;
        RECT 95.330 74.405 96.980 74.575 ;
        RECT 96.810 74.335 96.980 74.405 ;
        RECT 96.810 74.165 97.455 74.335 ;
        RECT 94.070 73.945 94.240 74.050 ;
        RECT 97.285 74.135 97.455 74.165 ;
        RECT 97.285 73.965 102.475 74.135 ;
        RECT 94.070 73.775 96.875 73.945 ;
        RECT 79.525 73.060 80.145 73.390 ;
        RECT 90.890 72.545 91.890 73.545 ;
        RECT 96.705 73.505 96.875 73.775 ;
        RECT 93.130 73.295 96.515 73.465 ;
        RECT 96.705 73.335 102.475 73.505 ;
        RECT 93.130 73.230 93.300 73.295 ;
        RECT 92.770 73.060 93.300 73.230 ;
        RECT 93.925 72.770 95.790 72.940 ;
        RECT 89.570 72.330 90.100 72.415 ;
        RECT 89.570 72.160 90.360 72.330 ;
        RECT 51.105 71.930 52.170 72.025 ;
        RECT 51.105 71.760 52.270 71.930 ;
        RECT 90.190 71.760 90.360 72.160 ;
        RECT 91.540 72.220 91.710 72.545 ;
        RECT 93.925 72.220 94.095 72.770 ;
        RECT 91.540 72.050 94.095 72.220 ;
        RECT 95.620 72.245 95.790 72.770 ;
        RECT 96.345 72.875 96.515 73.295 ;
        RECT 96.345 72.705 102.475 72.875 ;
        RECT 95.620 72.075 102.475 72.245 ;
        RECT 91.180 71.760 93.455 71.785 ;
        RECT 51.105 71.695 52.170 71.760 ;
        RECT 51.105 67.445 51.435 71.695 ;
        RECT 51.870 70.975 52.040 71.695 ;
        RECT 90.190 71.615 93.455 71.760 ;
        RECT 90.190 71.590 91.350 71.615 ;
        RECT 93.285 71.445 102.475 71.615 ;
        RECT 87.675 70.985 88.675 71.405 ;
        RECT 51.860 70.805 57.630 70.975 ;
        RECT 87.675 70.815 102.475 70.985 ;
        RECT 87.675 70.405 88.675 70.815 ;
        RECT 97.725 70.325 102.475 70.355 ;
        RECT 96.200 70.185 102.475 70.325 ;
        RECT 96.200 70.155 97.955 70.185 ;
        RECT 96.200 70.055 96.370 70.155 ;
        RECT 89.570 69.885 96.370 70.055 ;
        RECT 96.765 69.725 97.905 69.740 ;
        RECT 75.660 69.430 76.190 69.605 ;
        RECT 96.765 69.570 102.475 69.725 ;
        RECT 96.765 69.520 96.935 69.570 ;
        RECT 97.725 69.555 102.475 69.570 ;
        RECT 75.660 69.260 83.670 69.430 ;
        RECT 75.660 69.075 76.190 69.260 ;
        RECT 63.915 68.960 64.645 68.965 ;
        RECT 63.735 68.950 64.645 68.960 ;
        RECT 58.270 68.285 58.800 68.815 ;
        RECT 63.735 68.795 71.315 68.950 ;
        RECT 63.735 68.790 64.265 68.795 ;
        RECT 64.525 68.780 71.315 68.795 ;
        RECT 61.585 67.870 71.315 68.040 ;
        RECT 51.860 67.675 57.630 67.695 ;
        RECT 51.850 67.525 57.630 67.675 ;
        RECT 51.850 67.060 52.020 67.525 ;
        RECT 51.390 66.060 52.390 67.060 ;
        RECT 61.585 66.220 61.755 67.870 ;
        RECT 63.915 67.140 64.775 67.145 ;
        RECT 63.735 67.130 64.775 67.140 ;
        RECT 63.735 66.975 71.315 67.130 ;
        RECT 63.735 66.970 64.265 66.975 ;
        RECT 64.525 66.960 71.315 66.975 ;
        RECT 61.585 66.050 71.315 66.220 ;
        RECT 51.105 65.390 52.170 65.420 ;
        RECT 51.105 65.220 52.270 65.390 ;
        RECT 51.105 65.090 52.170 65.220 ;
        RECT 51.105 60.755 51.435 65.090 ;
        RECT 51.860 64.285 52.030 65.090 ;
        RECT 61.585 64.400 61.755 66.050 ;
        RECT 63.915 65.320 64.755 65.325 ;
        RECT 63.735 65.310 64.755 65.320 ;
        RECT 63.735 65.155 71.315 65.310 ;
        RECT 63.735 65.150 64.265 65.155 ;
        RECT 64.525 65.140 71.315 65.155 ;
        RECT 51.860 64.115 57.630 64.285 ;
        RECT 61.585 64.230 71.315 64.400 ;
        RECT 58.290 62.950 58.820 63.480 ;
        RECT 61.585 62.580 61.755 64.230 ;
        RECT 63.745 63.490 64.645 63.505 ;
        RECT 63.745 63.335 71.315 63.490 ;
        RECT 64.525 63.320 71.315 63.335 ;
        RECT 61.585 62.410 71.315 62.580 ;
        RECT 51.860 60.985 57.630 61.005 ;
        RECT 51.850 60.835 57.630 60.985 ;
        RECT 51.850 60.370 52.020 60.835 ;
        RECT 61.585 60.760 61.755 62.410 ;
        RECT 63.745 61.670 64.275 61.680 ;
        RECT 63.745 61.510 71.315 61.670 ;
        RECT 63.925 61.500 71.315 61.510 ;
        RECT 61.585 60.590 71.315 60.760 ;
        RECT 51.390 59.370 52.390 60.370 ;
        RECT 61.585 58.940 61.755 60.590 ;
        RECT 63.925 59.855 64.790 59.865 ;
        RECT 63.745 59.850 64.790 59.855 ;
        RECT 63.745 59.695 71.315 59.850 ;
        RECT 63.745 59.685 64.275 59.695 ;
        RECT 64.525 59.680 71.315 59.695 ;
        RECT 61.585 58.770 71.315 58.940 ;
        RECT 51.105 58.695 52.170 58.765 ;
        RECT 51.105 58.525 52.270 58.695 ;
        RECT 51.105 58.435 52.170 58.525 ;
        RECT 51.105 54.065 51.435 58.435 ;
        RECT 51.865 57.595 52.035 58.435 ;
        RECT 61.585 57.930 61.755 58.770 ;
        RECT 63.735 58.030 64.780 58.045 ;
        RECT 62.155 57.930 62.425 58.015 ;
        RECT 61.585 57.760 62.425 57.930 ;
        RECT 63.735 57.875 71.315 58.030 ;
        RECT 64.525 57.860 71.315 57.875 ;
        RECT 51.860 57.425 57.630 57.595 ;
        RECT 61.585 57.120 61.755 57.760 ;
        RECT 62.155 57.685 62.425 57.760 ;
        RECT 61.585 56.950 71.315 57.120 ;
        RECT 61.585 56.220 61.755 56.950 ;
        RECT 64.010 56.225 64.205 56.340 ;
        RECT 64.010 56.220 64.740 56.225 ;
        RECT 61.440 56.050 61.970 56.220 ;
        RECT 63.745 56.210 64.740 56.220 ;
        RECT 63.745 56.055 71.315 56.210 ;
        RECT 71.730 56.195 72.060 69.030 ;
        RECT 74.460 67.980 83.670 68.150 ;
        RECT 74.510 65.590 74.680 67.980 ;
        RECT 75.660 66.870 76.190 67.090 ;
        RECT 75.660 66.700 83.670 66.870 ;
        RECT 75.660 66.560 76.190 66.700 ;
        RECT 74.510 65.420 83.670 65.590 ;
        RECT 74.510 63.030 74.680 65.420 ;
        RECT 75.660 64.310 76.190 64.485 ;
        RECT 75.660 64.140 83.670 64.310 ;
        RECT 75.660 63.955 76.190 64.140 ;
        RECT 74.510 62.860 83.670 63.030 ;
        RECT 74.510 60.470 74.680 62.860 ;
        RECT 75.660 61.750 76.190 61.955 ;
        RECT 75.660 61.580 83.670 61.750 ;
        RECT 75.660 61.425 76.190 61.580 ;
        RECT 74.510 60.300 83.670 60.470 ;
        RECT 74.510 57.910 74.680 60.300 ;
        RECT 75.660 59.190 76.190 59.310 ;
        RECT 75.660 59.020 83.670 59.190 ;
        RECT 75.660 58.780 76.190 59.020 ;
        RECT 74.510 57.740 83.670 57.910 ;
        RECT 74.510 57.330 74.680 57.740 ;
        RECT 74.510 57.180 74.785 57.330 ;
        RECT 74.515 57.000 74.785 57.180 ;
        RECT 63.745 56.050 64.275 56.055 ;
        RECT 64.525 56.040 71.315 56.055 ;
        RECT 71.710 55.960 72.060 56.195 ;
        RECT 74.540 56.165 74.710 57.000 ;
        RECT 75.660 56.630 76.190 56.835 ;
        RECT 75.660 56.460 83.670 56.630 ;
        RECT 75.660 56.305 76.190 56.460 ;
        RECT 84.085 56.380 84.415 69.510 ;
        RECT 90.625 69.350 96.935 69.520 ;
        RECT 90.625 69.005 90.795 69.350 ;
        RECT 97.725 69.075 102.475 69.095 ;
        RECT 97.225 69.035 102.475 69.075 ;
        RECT 90.210 68.005 91.210 69.005 ;
        RECT 92.350 68.925 102.475 69.035 ;
        RECT 92.350 68.905 97.895 68.925 ;
        RECT 92.350 68.865 97.395 68.905 ;
        RECT 92.350 68.590 92.520 68.865 ;
        RECT 91.905 68.420 92.520 68.590 ;
        RECT 93.005 68.295 102.475 68.465 ;
        RECT 93.005 67.580 93.175 68.295 ;
        RECT 94.470 67.665 102.475 67.835 ;
        RECT 92.285 66.580 93.285 67.580 ;
        RECT 94.470 67.070 94.640 67.665 ;
        RECT 94.010 66.900 94.640 67.070 ;
        RECT 94.190 66.860 94.640 66.900 ;
        RECT 95.180 67.035 102.475 67.205 ;
        RECT 95.180 66.165 95.350 67.035 ;
        RECT 93.160 65.995 95.350 66.165 ;
        RECT 95.790 66.405 102.475 66.575 ;
        RECT 93.160 65.635 93.330 65.995 ;
        RECT 92.285 65.050 93.330 65.635 ;
        RECT 95.790 65.315 95.960 66.405 ;
        RECT 94.395 65.245 95.960 65.315 ;
        RECT 94.215 65.145 95.960 65.245 ;
        RECT 96.410 65.775 102.475 65.945 ;
        RECT 94.215 65.075 94.745 65.145 ;
        RECT 92.285 64.635 93.285 65.050 ;
        RECT 96.410 64.760 96.580 65.775 ;
        RECT 102.910 65.490 103.240 76.735 ;
        RECT 112.920 75.395 113.920 76.370 ;
        RECT 114.585 76.210 115.115 76.235 ;
        RECT 114.585 76.065 115.200 76.210 ;
        RECT 114.955 76.040 115.200 76.065 ;
        RECT 112.920 75.370 114.760 75.395 ;
        RECT 113.495 75.225 114.760 75.370 ;
        RECT 111.890 73.805 112.890 74.805 ;
        RECT 114.590 74.735 114.760 75.225 ;
        RECT 115.030 75.150 115.200 76.040 ;
        RECT 115.550 75.770 115.720 77.095 ;
        RECT 116.695 76.410 116.865 77.315 ;
        RECT 116.380 76.240 121.130 76.410 ;
        RECT 116.380 75.770 121.130 75.780 ;
        RECT 115.550 75.610 121.130 75.770 ;
        RECT 115.550 75.600 116.520 75.610 ;
        RECT 115.030 74.980 121.130 75.150 ;
        RECT 114.590 74.565 116.090 74.735 ;
        RECT 113.535 74.395 114.150 74.565 ;
        RECT 113.980 74.330 114.150 74.395 ;
        RECT 115.920 74.520 116.090 74.565 ;
        RECT 115.920 74.350 121.130 74.520 ;
        RECT 113.980 74.160 115.630 74.330 ;
        RECT 115.460 74.090 115.630 74.160 ;
        RECT 115.460 73.920 116.105 74.090 ;
        RECT 112.720 73.700 112.890 73.805 ;
        RECT 115.935 73.890 116.105 73.920 ;
        RECT 115.935 73.720 121.130 73.890 ;
        RECT 112.720 73.530 115.525 73.700 ;
        RECT 109.540 72.300 110.540 73.300 ;
        RECT 115.355 73.260 115.525 73.530 ;
        RECT 111.780 73.050 115.165 73.220 ;
        RECT 115.355 73.090 121.130 73.260 ;
        RECT 111.780 72.985 111.950 73.050 ;
        RECT 111.420 72.815 111.950 72.985 ;
        RECT 112.575 72.525 114.440 72.695 ;
        RECT 108.220 72.085 108.750 72.170 ;
        RECT 108.220 71.915 109.010 72.085 ;
        RECT 108.840 71.515 109.010 71.915 ;
        RECT 110.190 71.975 110.360 72.300 ;
        RECT 112.575 71.975 112.745 72.525 ;
        RECT 110.190 71.805 112.745 71.975 ;
        RECT 114.270 72.000 114.440 72.525 ;
        RECT 114.995 72.630 115.165 73.050 ;
        RECT 114.995 72.460 121.130 72.630 ;
        RECT 114.270 71.830 121.130 72.000 ;
        RECT 109.830 71.515 112.105 71.540 ;
        RECT 108.840 71.370 112.105 71.515 ;
        RECT 108.840 71.345 110.000 71.370 ;
        RECT 111.935 71.200 121.130 71.370 ;
        RECT 106.325 70.740 107.325 71.175 ;
        RECT 121.565 71.045 121.895 76.490 ;
        RECT 106.325 70.570 121.130 70.740 ;
        RECT 106.325 70.175 107.325 70.570 ;
        RECT 121.565 70.345 122.730 71.045 ;
        RECT 116.380 70.080 121.130 70.110 ;
        RECT 114.850 69.940 121.130 70.080 ;
        RECT 114.850 69.910 116.605 69.940 ;
        RECT 114.850 69.810 115.020 69.910 ;
        RECT 108.220 69.640 115.020 69.810 ;
        RECT 115.415 69.480 116.555 69.495 ;
        RECT 115.415 69.325 121.130 69.480 ;
        RECT 115.415 69.275 115.585 69.325 ;
        RECT 116.380 69.310 121.130 69.325 ;
        RECT 109.275 69.105 115.585 69.275 ;
        RECT 109.275 68.760 109.445 69.105 ;
        RECT 116.380 68.830 121.130 68.850 ;
        RECT 115.875 68.790 121.130 68.830 ;
        RECT 108.860 67.760 109.860 68.760 ;
        RECT 111.000 68.680 121.130 68.790 ;
        RECT 111.000 68.660 116.545 68.680 ;
        RECT 111.000 68.620 116.045 68.660 ;
        RECT 111.000 68.345 111.170 68.620 ;
        RECT 110.555 68.175 111.170 68.345 ;
        RECT 111.655 68.050 121.130 68.220 ;
        RECT 111.655 67.335 111.825 68.050 ;
        RECT 113.120 67.420 121.130 67.590 ;
        RECT 110.935 66.335 111.935 67.335 ;
        RECT 113.120 66.825 113.290 67.420 ;
        RECT 112.660 66.655 113.290 66.825 ;
        RECT 112.840 66.615 113.290 66.655 ;
        RECT 113.830 66.790 121.130 66.960 ;
        RECT 113.830 65.920 114.000 66.790 ;
        RECT 111.810 65.750 114.000 65.920 ;
        RECT 114.440 66.160 121.130 66.330 ;
        RECT 104.100 65.490 104.630 65.605 ;
        RECT 95.350 64.590 96.580 64.760 ;
        RECT 96.900 65.145 102.475 65.315 ;
        RECT 102.910 65.190 104.630 65.490 ;
        RECT 111.810 65.390 111.980 65.750 ;
        RECT 95.350 64.095 95.520 64.590 ;
        RECT 94.555 63.095 95.555 64.095 ;
        RECT 96.900 63.820 97.070 65.145 ;
        RECT 97.725 64.515 102.475 64.685 ;
        RECT 98.125 64.095 98.295 64.515 ;
        RECT 102.910 64.435 103.240 65.190 ;
        RECT 104.100 65.075 104.630 65.190 ;
        RECT 110.935 64.805 111.980 65.390 ;
        RECT 114.440 65.070 114.610 66.160 ;
        RECT 113.045 65.000 114.610 65.070 ;
        RECT 112.865 64.900 114.610 65.000 ;
        RECT 115.060 65.530 121.130 65.700 ;
        RECT 112.865 64.830 113.395 64.900 ;
        RECT 110.935 64.390 111.935 64.805 ;
        RECT 115.060 64.515 115.230 65.530 ;
        RECT 114.000 64.345 115.230 64.515 ;
        RECT 115.550 64.900 121.130 65.070 ;
        RECT 96.475 63.785 97.070 63.820 ;
        RECT 96.295 63.650 97.070 63.785 ;
        RECT 96.295 63.615 96.825 63.650 ;
        RECT 97.710 63.095 98.710 64.095 ;
        RECT 114.000 63.850 114.170 64.345 ;
        RECT 113.205 62.850 114.205 63.850 ;
        RECT 115.550 63.575 115.720 64.900 ;
        RECT 116.380 64.270 121.130 64.440 ;
        RECT 116.775 63.850 116.945 64.270 ;
        RECT 121.565 64.190 121.895 70.345 ;
        RECT 115.125 63.540 115.720 63.575 ;
        RECT 114.945 63.405 115.720 63.540 ;
        RECT 114.945 63.370 115.475 63.405 ;
        RECT 116.360 62.850 117.360 63.850 ;
        RECT 107.210 57.740 107.875 57.910 ;
        RECT 71.710 55.695 72.010 55.960 ;
        RECT 71.710 55.395 72.255 55.695 ;
        RECT 74.335 55.635 74.865 56.165 ;
        RECT 58.270 54.465 58.800 54.995 ;
        RECT 51.850 54.315 52.020 54.320 ;
        RECT 51.850 54.145 57.630 54.315 ;
        RECT 71.955 54.150 72.255 55.395 ;
        RECT 84.090 54.320 84.390 56.380 ;
        RECT 106.310 56.335 107.310 56.805 ;
        RECT 107.705 56.795 107.875 57.740 ;
        RECT 108.560 57.215 109.560 58.215 ;
        RECT 110.215 57.740 110.995 57.910 ;
        RECT 109.295 57.005 109.465 57.215 ;
        RECT 109.295 56.835 110.500 57.005 ;
        RECT 107.705 56.625 108.965 56.795 ;
        RECT 108.795 56.370 108.965 56.625 ;
        RECT 106.310 56.165 108.450 56.335 ;
        RECT 108.795 56.200 110.005 56.370 ;
        RECT 106.310 55.805 107.310 56.165 ;
        RECT 108.280 55.810 108.450 56.165 ;
        RECT 108.280 55.640 109.480 55.810 ;
        RECT 109.310 55.190 109.480 55.640 ;
        RECT 109.835 55.700 110.005 56.200 ;
        RECT 110.330 56.215 110.500 56.835 ;
        RECT 110.825 56.735 110.995 57.740 ;
        RECT 111.560 57.800 112.560 58.215 ;
        RECT 111.560 57.215 112.630 57.800 ;
        RECT 110.825 56.565 112.160 56.735 ;
        RECT 110.330 56.045 111.680 56.215 ;
        RECT 109.835 55.530 111.220 55.700 ;
        RECT 84.090 54.150 84.420 54.320 ;
        RECT 51.850 53.705 52.020 54.145 ;
        RECT 51.390 52.705 52.390 53.705 ;
        RECT 71.840 53.620 72.370 54.150 ;
        RECT 83.995 53.620 84.525 54.150 ;
        RECT 105.975 54.130 106.975 55.130 ;
        RECT 109.310 55.020 110.705 55.190 ;
        RECT 107.765 54.665 108.830 54.835 ;
        RECT 108.660 54.595 108.830 54.665 ;
        RECT 108.660 54.425 110.205 54.595 ;
        RECT 106.645 53.785 106.815 54.130 ;
        RECT 51.105 51.635 52.195 51.965 ;
        RECT 60.020 51.920 60.910 52.810 ;
        RECT 64.150 52.255 64.880 52.260 ;
        RECT 63.970 52.245 64.880 52.255 ;
        RECT 63.970 52.090 71.570 52.245 ;
        RECT 63.970 52.085 64.500 52.090 ;
        RECT 64.780 52.075 71.570 52.090 ;
        RECT 51.105 47.425 51.435 51.635 ;
        RECT 51.665 51.595 52.195 51.635 ;
        RECT 51.860 50.955 52.030 51.595 ;
        RECT 61.405 51.335 62.405 51.815 ;
        RECT 61.405 51.165 71.570 51.335 ;
        RECT 51.860 50.785 57.630 50.955 ;
        RECT 61.405 50.815 62.405 51.165 ;
        RECT 64.150 50.435 65.010 50.440 ;
        RECT 63.970 50.425 65.010 50.435 ;
        RECT 63.970 50.270 71.570 50.425 ;
        RECT 63.970 50.265 64.500 50.270 ;
        RECT 64.780 50.255 71.570 50.270 ;
        RECT 61.405 49.515 62.405 49.930 ;
        RECT 58.290 48.895 58.820 49.425 ;
        RECT 61.405 49.345 71.570 49.515 ;
        RECT 61.405 48.930 62.405 49.345 ;
        RECT 64.150 48.615 64.990 48.620 ;
        RECT 63.970 48.605 64.990 48.615 ;
        RECT 63.970 48.450 71.570 48.605 ;
        RECT 63.970 48.445 64.500 48.450 ;
        RECT 64.780 48.435 71.570 48.450 ;
        RECT 61.405 47.695 62.405 48.105 ;
        RECT 51.850 47.675 52.020 47.695 ;
        RECT 51.850 47.505 57.630 47.675 ;
        RECT 61.405 47.525 71.570 47.695 ;
        RECT 51.850 47.080 52.020 47.505 ;
        RECT 61.405 47.105 62.405 47.525 ;
        RECT 37.260 45.160 38.510 46.410 ;
        RECT 51.390 46.080 52.390 47.080 ;
        RECT 63.980 46.780 64.510 46.795 ;
        RECT 64.780 46.780 71.570 46.785 ;
        RECT 63.980 46.625 71.570 46.780 ;
        RECT 64.160 46.615 71.570 46.625 ;
        RECT 64.160 46.610 64.880 46.615 ;
        RECT 61.405 45.875 62.405 46.230 ;
        RECT 61.405 45.705 71.570 45.875 ;
        RECT 43.830 45.295 44.360 45.465 ;
        RECT 37.635 44.835 37.935 45.160 ;
        RECT 37.635 41.225 37.965 44.835 ;
        RECT 44.005 44.755 44.175 45.295 ;
        RECT 48.405 45.290 48.935 45.460 ;
        RECT 38.440 44.585 44.210 44.755 ;
        RECT 44.005 44.575 44.175 44.585 ;
        RECT 47.760 43.435 48.090 44.835 ;
        RECT 48.580 44.755 48.750 45.290 ;
        RECT 61.405 45.230 62.405 45.705 ;
        RECT 63.980 44.960 64.510 44.975 ;
        RECT 64.780 44.960 71.570 44.965 ;
        RECT 63.980 44.805 71.570 44.960 ;
        RECT 64.160 44.795 71.570 44.805 ;
        RECT 64.160 44.790 64.930 44.795 ;
        RECT 48.565 44.585 54.335 44.755 ;
        RECT 48.580 44.570 48.750 44.585 ;
        RECT 47.005 43.320 48.090 43.435 ;
        RECT 61.405 44.055 62.405 44.410 ;
        RECT 61.405 43.885 71.570 44.055 ;
        RECT 61.405 43.410 62.405 43.885 ;
        RECT 44.990 42.735 45.520 43.265 ;
        RECT 46.905 43.150 48.090 43.320 ;
        RECT 64.160 43.150 65.025 43.160 ;
        RECT 47.005 43.105 48.090 43.150 ;
        RECT 38.440 41.305 44.210 41.475 ;
        RECT 39.775 40.850 39.945 41.305 ;
        RECT 47.760 41.225 48.090 43.105 ;
        RECT 63.980 43.145 65.025 43.150 ;
        RECT 63.980 42.990 71.570 43.145 ;
        RECT 63.980 42.980 64.510 42.990 ;
        RECT 64.780 42.975 71.570 42.990 ;
        RECT 55.050 42.320 55.580 42.850 ;
        RECT 61.405 42.235 62.405 42.670 ;
        RECT 61.405 42.065 71.570 42.235 ;
        RECT 61.405 41.670 62.405 42.065 ;
        RECT 48.565 41.305 54.335 41.475 ;
        RECT 63.970 41.325 65.015 41.340 ;
        RECT 48.585 40.860 48.755 41.305 ;
        RECT 63.970 41.170 71.570 41.325 ;
        RECT 64.780 41.155 71.570 41.170 ;
        RECT 39.315 39.850 40.315 40.850 ;
        RECT 48.125 39.860 49.125 40.860 ;
        RECT 61.405 40.415 62.405 40.835 ;
        RECT 61.405 40.245 71.570 40.415 ;
        RECT 61.405 39.835 62.405 40.245 ;
        RECT 37.260 38.430 38.510 39.680 ;
        RECT 64.245 39.520 64.440 39.635 ;
        RECT 64.245 39.515 64.975 39.520 ;
        RECT 63.980 39.505 64.975 39.515 ;
        RECT 63.980 39.350 71.570 39.505 ;
        RECT 63.980 39.345 64.510 39.350 ;
        RECT 64.780 39.335 71.570 39.350 ;
        RECT 71.985 39.255 72.315 53.620 ;
        RECT 74.660 51.785 75.270 52.455 ;
        RECT 75.660 51.780 76.190 51.960 ;
        RECT 84.090 51.865 84.420 53.620 ;
        RECT 106.645 53.615 109.610 53.785 ;
        RECT 106.905 52.660 108.760 52.665 ;
        RECT 106.725 52.495 108.760 52.660 ;
        RECT 106.725 52.490 107.255 52.495 ;
        RECT 76.900 51.780 83.690 51.785 ;
        RECT 75.660 51.615 83.690 51.780 ;
        RECT 84.090 51.655 84.435 51.865 ;
        RECT 75.660 51.610 77.080 51.615 ;
        RECT 75.660 51.430 76.190 51.610 ;
        RECT 72.940 50.500 73.940 50.930 ;
        RECT 76.900 50.500 83.690 50.505 ;
        RECT 72.940 50.335 83.690 50.500 ;
        RECT 72.940 50.330 77.075 50.335 ;
        RECT 72.940 49.930 73.940 50.330 ;
        RECT 75.585 49.220 76.115 49.395 ;
        RECT 76.900 49.220 83.690 49.225 ;
        RECT 75.585 49.055 83.690 49.220 ;
        RECT 75.585 49.050 76.970 49.055 ;
        RECT 75.585 48.865 76.115 49.050 ;
        RECT 72.880 47.940 73.880 48.360 ;
        RECT 76.900 47.940 83.690 47.945 ;
        RECT 72.880 47.775 83.690 47.940 ;
        RECT 72.880 47.770 76.970 47.775 ;
        RECT 72.880 47.360 73.880 47.770 ;
        RECT 75.580 46.660 76.110 46.840 ;
        RECT 76.900 46.660 83.690 46.665 ;
        RECT 75.580 46.495 83.690 46.660 ;
        RECT 75.580 46.490 76.970 46.495 ;
        RECT 75.580 46.310 76.110 46.490 ;
        RECT 72.990 45.380 73.990 45.855 ;
        RECT 76.900 45.380 83.690 45.385 ;
        RECT 72.990 45.215 83.690 45.380 ;
        RECT 72.990 45.210 76.970 45.215 ;
        RECT 72.990 44.855 73.990 45.210 ;
        RECT 75.620 44.100 76.150 44.275 ;
        RECT 76.900 44.100 83.690 44.105 ;
        RECT 75.620 43.935 83.690 44.100 ;
        RECT 75.620 43.930 76.970 43.935 ;
        RECT 75.620 43.745 76.150 43.930 ;
        RECT 72.990 42.820 73.990 43.245 ;
        RECT 76.900 42.820 83.690 42.825 ;
        RECT 72.990 42.655 83.690 42.820 ;
        RECT 72.990 42.650 76.970 42.655 ;
        RECT 72.990 42.245 73.990 42.650 ;
        RECT 75.595 41.540 76.125 41.715 ;
        RECT 76.900 41.540 83.690 41.545 ;
        RECT 75.595 41.375 83.690 41.540 ;
        RECT 75.595 41.370 76.970 41.375 ;
        RECT 75.595 41.185 76.125 41.370 ;
        RECT 72.990 40.260 73.990 40.760 ;
        RECT 76.900 40.260 83.690 40.265 ;
        RECT 72.990 40.095 83.690 40.260 ;
        RECT 72.990 40.090 76.970 40.095 ;
        RECT 72.990 39.760 73.990 40.090 ;
        RECT 43.850 38.635 44.380 38.805 ;
        RECT 48.405 38.660 48.935 38.830 ;
        RECT 76.900 38.815 83.690 38.985 ;
        RECT 37.640 38.140 37.960 38.430 ;
        RECT 37.635 34.530 37.965 38.140 ;
        RECT 44.025 38.060 44.195 38.635 ;
        RECT 38.440 37.890 44.210 38.060 ;
        RECT 44.960 36.030 45.490 36.560 ;
        RECT 47.760 36.390 48.090 38.140 ;
        RECT 48.580 38.060 48.750 38.660 ;
        RECT 76.070 38.110 76.600 38.290 ;
        RECT 77.660 38.110 77.830 38.815 ;
        RECT 84.105 38.735 84.435 51.655 ;
        RECT 108.590 51.710 108.760 52.495 ;
        RECT 109.440 52.340 109.610 53.615 ;
        RECT 110.035 52.970 110.205 54.425 ;
        RECT 110.535 53.600 110.705 55.020 ;
        RECT 111.050 54.230 111.220 55.530 ;
        RECT 111.510 54.860 111.680 56.045 ;
        RECT 111.990 55.490 112.160 56.565 ;
        RECT 112.460 56.120 112.630 57.215 ;
        RECT 114.100 56.750 114.800 57.910 ;
        RECT 113.545 56.580 120.335 56.750 ;
        RECT 112.460 55.950 120.335 56.120 ;
        RECT 111.990 55.320 120.335 55.490 ;
        RECT 111.510 54.690 120.335 54.860 ;
        RECT 111.050 54.060 120.335 54.230 ;
        RECT 110.535 53.430 120.335 53.600 ;
        RECT 110.035 52.800 120.335 52.970 ;
        RECT 109.440 52.170 120.335 52.340 ;
        RECT 120.750 51.715 121.080 56.830 ;
        RECT 108.590 51.540 120.335 51.710 ;
        RECT 105.975 51.080 106.975 51.510 ;
        RECT 105.975 50.910 120.335 51.080 ;
        RECT 120.750 51.015 122.455 51.715 ;
        RECT 105.975 50.510 106.975 50.910 ;
        RECT 108.430 50.280 120.335 50.450 ;
        RECT 108.430 49.385 108.600 50.280 ;
        RECT 106.905 49.380 108.600 49.385 ;
        RECT 106.725 49.215 108.600 49.380 ;
        RECT 109.320 49.820 113.710 49.830 ;
        RECT 109.320 49.660 120.335 49.820 ;
        RECT 106.725 49.210 107.255 49.215 ;
        RECT 109.320 48.520 109.490 49.660 ;
        RECT 113.545 49.650 120.335 49.660 ;
        RECT 108.525 48.350 109.490 48.520 ;
        RECT 109.930 49.020 120.335 49.190 ;
        RECT 108.525 48.265 108.695 48.350 ;
        RECT 106.390 48.095 108.695 48.265 ;
        RECT 106.390 47.760 106.560 48.095 ;
        RECT 109.930 47.845 110.100 49.020 ;
        RECT 105.975 46.760 106.975 47.760 ;
        RECT 109.135 47.675 110.100 47.845 ;
        RECT 110.455 48.390 120.335 48.560 ;
        RECT 109.135 47.340 109.305 47.675 ;
        RECT 107.765 47.170 109.305 47.340 ;
        RECT 110.455 47.225 110.625 48.390 ;
        RECT 109.675 47.055 110.625 47.225 ;
        RECT 111.040 47.760 120.335 47.930 ;
        RECT 109.675 46.225 109.845 47.055 ;
        RECT 111.040 46.645 111.210 47.760 ;
        RECT 106.650 45.670 107.650 46.155 ;
        RECT 108.685 46.055 109.845 46.225 ;
        RECT 110.215 46.475 111.210 46.645 ;
        RECT 111.530 47.130 120.335 47.300 ;
        RECT 108.685 45.670 108.855 46.055 ;
        RECT 106.650 45.500 108.855 45.670 ;
        RECT 110.215 45.645 110.385 46.475 ;
        RECT 111.530 46.035 111.700 47.130 ;
        RECT 106.650 45.155 107.650 45.500 ;
        RECT 109.350 45.475 110.385 45.645 ;
        RECT 110.735 45.865 111.700 46.035 ;
        RECT 112.090 46.500 120.335 46.670 ;
        RECT 109.350 45.210 109.520 45.475 ;
        RECT 108.260 45.040 109.520 45.210 ;
        RECT 110.735 45.160 110.905 45.865 ;
        RECT 112.090 45.395 112.260 46.500 ;
        RECT 108.260 44.210 108.430 45.040 ;
        RECT 109.900 44.990 110.905 45.160 ;
        RECT 111.245 45.225 112.260 45.395 ;
        RECT 112.750 45.870 120.335 46.040 ;
        RECT 109.900 44.665 110.070 44.990 ;
        RECT 107.765 44.040 108.430 44.210 ;
        RECT 107.945 44.030 108.430 44.040 ;
        RECT 109.060 44.080 110.070 44.665 ;
        RECT 111.245 44.210 111.415 45.225 ;
        RECT 112.750 44.705 112.920 45.870 ;
        RECT 113.545 45.240 120.335 45.410 ;
        RECT 114.355 45.235 114.535 45.240 ;
        RECT 110.845 44.185 111.415 44.210 ;
        RECT 109.060 43.665 110.060 44.080 ;
        RECT 110.665 44.040 111.415 44.185 ;
        RECT 111.790 44.135 112.920 44.705 ;
        RECT 114.365 44.440 114.535 45.235 ;
        RECT 120.750 45.160 121.080 51.015 ;
        RECT 114.185 44.270 114.715 44.440 ;
        RECT 110.665 44.015 111.195 44.040 ;
        RECT 111.790 43.705 112.790 44.135 ;
        RECT 112.775 41.675 113.305 42.205 ;
        RECT 48.565 37.890 54.335 38.060 ;
        RECT 76.070 37.940 77.830 38.110 ;
        RECT 76.070 37.760 76.600 37.940 ;
        RECT 57.865 36.515 58.395 36.845 ;
        RECT 47.005 36.355 48.090 36.390 ;
        RECT 46.905 36.185 48.090 36.355 ;
        RECT 47.005 36.060 48.090 36.185 ;
        RECT 38.440 34.610 44.210 34.780 ;
        RECT 39.425 34.145 39.595 34.610 ;
        RECT 47.760 34.530 48.090 36.060 ;
        RECT 55.070 35.985 55.600 36.515 ;
        RECT 58.065 35.160 58.395 36.515 ;
        RECT 58.965 35.625 59.965 36.625 ;
        RECT 72.860 36.040 73.750 36.930 ;
        RECT 58.665 35.160 58.995 35.205 ;
        RECT 58.065 34.830 58.995 35.160 ;
        RECT 59.465 35.125 59.635 35.625 ;
        RECT 59.410 34.955 66.200 35.125 ;
        RECT 48.565 34.610 54.335 34.780 ;
        RECT 48.570 34.155 48.740 34.610 ;
        RECT 37.260 32.335 38.510 33.585 ;
        RECT 38.965 33.145 39.965 34.145 ;
        RECT 48.110 33.155 49.110 34.155 ;
        RECT 58.665 33.965 58.995 34.830 ;
        RECT 66.570 34.265 67.180 34.935 ;
        RECT 72.115 34.910 72.445 35.380 ;
        RECT 73.295 35.300 73.465 36.040 ;
        RECT 72.860 35.130 79.650 35.300 ;
        RECT 71.045 34.850 72.445 34.910 ;
        RECT 70.945 34.680 72.445 34.850 ;
        RECT 71.045 34.580 72.445 34.680 ;
        RECT 59.410 34.045 66.200 34.215 ;
        RECT 72.115 34.140 72.445 34.580 ;
        RECT 72.860 34.220 79.650 34.390 ;
        RECT 80.620 34.385 81.230 35.055 ;
        RECT 59.425 33.580 59.595 34.045 ;
        RECT 43.810 32.520 44.340 32.690 ;
        RECT 37.645 32.025 37.965 32.335 ;
        RECT 37.635 28.415 37.965 32.025 ;
        RECT 43.985 31.945 44.155 32.520 ;
        RECT 49.595 32.500 50.125 32.670 ;
        RECT 58.965 32.580 59.965 33.580 ;
        RECT 73.505 33.500 73.675 34.220 ;
        RECT 73.325 32.970 73.855 33.500 ;
        RECT 38.440 31.775 44.210 31.945 ;
        RECT 44.960 29.940 45.490 30.470 ;
        RECT 47.760 30.150 48.090 32.025 ;
        RECT 49.770 31.945 49.940 32.500 ;
        RECT 48.565 31.775 54.335 31.945 ;
        RECT 46.905 29.820 48.090 30.150 ;
        RECT 55.070 29.960 55.600 30.490 ;
        RECT 38.440 28.495 44.210 28.665 ;
        RECT 39.425 28.030 39.595 28.495 ;
        RECT 47.760 28.415 48.090 29.820 ;
        RECT 48.605 28.665 48.775 28.675 ;
        RECT 48.565 28.495 54.335 28.665 ;
        RECT 48.605 28.060 48.775 28.495 ;
        RECT 37.430 25.965 38.680 27.215 ;
        RECT 38.965 27.030 39.965 28.030 ;
        RECT 48.145 27.060 49.145 28.060 ;
        RECT 63.525 27.580 63.695 28.250 ;
        RECT 43.850 26.095 44.380 26.265 ;
        RECT 49.595 26.095 50.125 26.265 ;
        RECT 37.650 25.620 37.950 25.965 ;
        RECT 37.635 22.010 37.965 25.620 ;
        RECT 44.025 25.540 44.195 26.095 ;
        RECT 38.440 25.370 44.210 25.540 ;
        RECT 47.760 24.065 48.090 25.620 ;
        RECT 49.770 25.540 49.940 26.095 ;
        RECT 48.565 25.370 54.335 25.540 ;
        RECT 63.525 25.160 63.695 27.040 ;
        RECT 88.590 26.370 88.760 28.250 ;
        RECT 47.005 23.995 48.090 24.065 ;
        RECT 44.960 23.465 45.490 23.995 ;
        RECT 46.905 23.825 48.090 23.995 ;
        RECT 47.005 23.735 48.090 23.825 ;
        RECT 38.440 22.250 44.210 22.260 ;
        RECT 38.435 22.090 44.210 22.250 ;
        RECT 38.435 21.635 38.605 22.090 ;
        RECT 47.760 22.010 48.090 23.735 ;
        RECT 55.070 23.615 55.600 24.145 ;
        RECT 63.525 22.740 63.695 24.620 ;
        RECT 88.590 23.950 88.760 25.830 ;
        RECT 88.590 22.740 88.760 23.410 ;
        RECT 48.560 22.260 48.730 22.270 ;
        RECT 48.560 22.090 54.335 22.260 ;
        RECT 48.560 21.655 48.730 22.090 ;
        RECT 37.975 20.635 38.975 21.635 ;
        RECT 48.100 20.655 49.100 21.655 ;
      LAYER met1 ;
        RECT 59.880 219.530 88.945 219.600 ;
        RECT 59.835 218.630 88.945 219.530 ;
        RECT 59.880 218.600 88.945 218.630 ;
        RECT 59.880 216.055 60.880 218.600 ;
        RECT 87.945 216.055 88.945 218.600 ;
        RECT 37.435 214.665 43.110 216.055 ;
        RECT 10.695 213.665 43.110 214.665 ;
        RECT 37.435 210.415 43.110 213.665 ;
        RECT 56.055 210.555 66.055 216.055 ;
        RECT 83.795 210.645 93.795 216.055 ;
        RECT 119.930 215.945 124.435 216.055 ;
        RECT 119.930 214.945 128.520 215.945 ;
        RECT 95.510 213.765 114.440 214.465 ;
        RECT 37.435 209.715 54.265 210.415 ;
        RECT 37.435 185.960 43.110 209.715 ;
        RECT 51.480 208.395 52.180 209.715 ;
        RECT 51.480 207.695 52.235 208.395 ;
        RECT 51.500 205.350 52.200 207.695 ;
        RECT 58.750 207.490 59.340 208.140 ;
        RECT 53.275 205.770 53.865 206.420 ;
        RECT 51.500 204.650 54.255 205.350 ;
        RECT 51.500 203.495 52.200 204.650 ;
        RECT 51.500 202.795 52.235 203.495 ;
        RECT 58.895 203.485 59.195 207.490 ;
        RECT 62.435 206.000 63.135 210.555 ;
        RECT 63.850 206.700 64.440 207.350 ;
        RECT 91.345 206.000 92.045 210.645 ;
        RECT 92.935 206.700 93.525 207.350 ;
        RECT 62.310 204.990 63.260 206.000 ;
        RECT 91.220 204.990 92.170 206.000 ;
        RECT 58.750 202.835 59.340 203.485 ;
        RECT 63.670 202.895 64.260 203.545 ;
        RECT 92.935 202.915 93.525 203.565 ;
        RECT 51.520 198.920 52.220 202.795 ;
        RECT 53.235 200.960 53.825 201.610 ;
        RECT 51.520 198.220 54.180 198.920 ;
        RECT 51.520 196.260 52.275 198.220 ;
        RECT 58.895 197.090 59.195 202.835 ;
        RECT 95.510 202.605 96.210 213.765 ;
        RECT 98.735 213.175 99.325 213.350 ;
        RECT 93.690 202.590 96.210 202.605 ;
        RECT 63.675 201.785 64.255 202.425 ;
        RECT 64.890 201.905 96.210 202.590 ;
        RECT 96.650 212.875 99.325 213.175 ;
        RECT 96.650 205.980 96.950 212.875 ;
        RECT 98.735 212.700 99.325 212.875 ;
        RECT 104.360 211.895 104.960 213.765 ;
        RECT 107.015 213.095 107.605 213.350 ;
        RECT 104.345 211.245 104.960 211.895 ;
        RECT 97.370 210.080 97.970 210.720 ;
        RECT 102.800 206.910 103.390 207.560 ;
        RECT 98.735 205.980 99.325 206.155 ;
        RECT 96.650 205.680 99.325 205.980 ;
        RECT 64.890 201.890 94.390 201.905 ;
        RECT 64.890 201.820 65.590 201.890 ;
        RECT 58.750 196.440 59.340 197.090 ;
        RECT 51.520 193.995 52.220 196.260 ;
        RECT 53.290 195.015 53.880 195.190 ;
        RECT 58.895 195.015 59.195 196.440 ;
        RECT 53.290 194.715 59.195 195.015 ;
        RECT 53.290 194.540 53.880 194.715 ;
        RECT 51.520 193.295 54.235 193.995 ;
        RECT 51.520 192.270 52.220 193.295 ;
        RECT 51.520 191.570 52.235 192.270 ;
        RECT 58.895 192.045 59.195 194.715 ;
        RECT 58.750 191.395 59.340 192.045 ;
        RECT 53.290 190.195 53.880 190.370 ;
        RECT 58.895 190.195 59.195 191.395 ;
        RECT 53.290 189.895 59.195 190.195 ;
        RECT 53.290 189.720 53.880 189.895 ;
        RECT 53.435 187.440 53.735 189.720 ;
        RECT 53.225 186.800 53.805 187.440 ;
        RECT 37.435 185.910 47.055 185.960 ;
        RECT 37.435 185.260 55.635 185.910 ;
        RECT 37.435 181.230 43.110 185.260 ;
        RECT 44.340 184.000 45.040 185.260 ;
        RECT 46.355 185.210 55.635 185.260 ;
        RECT 53.610 183.125 54.200 183.775 ;
        RECT 52.600 181.775 53.190 181.950 ;
        RECT 53.755 181.775 54.055 183.125 ;
        RECT 54.215 181.775 54.795 181.940 ;
        RECT 52.600 181.475 54.795 181.775 ;
        RECT 52.600 181.300 53.190 181.475 ;
        RECT 37.435 180.530 47.000 181.230 ;
        RECT 37.435 176.655 43.110 180.530 ;
        RECT 44.330 179.545 45.030 180.530 ;
        RECT 53.755 179.320 54.055 181.475 ;
        RECT 54.215 181.300 54.795 181.475 ;
        RECT 53.610 178.670 54.200 179.320 ;
        RECT 52.600 177.260 53.190 177.435 ;
        RECT 53.755 177.260 54.055 178.670 ;
        RECT 52.600 176.960 54.055 177.260 ;
        RECT 52.600 176.785 53.190 176.960 ;
        RECT 37.435 176.640 46.890 176.655 ;
        RECT 37.435 175.990 47.000 176.640 ;
        RECT 37.435 175.955 46.890 175.990 ;
        RECT 37.435 171.115 43.110 175.955 ;
        RECT 44.330 174.945 45.030 175.955 ;
        RECT 53.755 174.625 54.055 176.960 ;
        RECT 54.935 175.545 55.635 185.210 ;
        RECT 56.400 184.115 56.980 184.290 ;
        RECT 63.815 184.115 64.115 201.785 ;
        RECT 83.070 200.290 83.770 201.890 ;
        RECT 81.300 199.590 83.770 200.290 ;
        RECT 75.990 197.495 76.570 198.135 ;
        RECT 76.150 197.105 76.450 197.495 ;
        RECT 76.015 196.455 76.605 197.105 ;
        RECT 76.150 194.035 76.450 196.455 ;
        RECT 77.460 194.035 78.050 194.210 ;
        RECT 76.150 193.735 78.050 194.035 ;
        RECT 76.150 189.830 76.450 193.735 ;
        RECT 77.460 193.560 78.050 193.735 ;
        RECT 83.070 193.185 83.770 199.590 ;
        RECT 81.300 192.485 83.770 193.185 ;
        RECT 83.070 191.385 83.770 192.485 ;
        RECT 96.650 199.005 96.950 205.680 ;
        RECT 98.735 205.505 99.325 205.680 ;
        RECT 97.370 202.905 97.970 203.545 ;
        RECT 102.885 199.845 103.475 200.495 ;
        RECT 98.735 199.005 99.325 199.180 ;
        RECT 96.650 198.705 99.325 199.005 ;
        RECT 96.650 191.995 96.950 198.705 ;
        RECT 98.735 198.530 99.325 198.705 ;
        RECT 97.370 195.955 97.970 196.595 ;
        RECT 102.885 192.965 103.475 193.615 ;
        RECT 98.735 191.995 99.325 192.205 ;
        RECT 96.650 191.695 99.325 191.995 ;
        RECT 75.995 189.180 76.585 189.830 ;
        RECT 76.140 187.205 76.440 189.180 ;
        RECT 95.600 188.880 96.200 189.520 ;
        RECT 77.460 187.205 78.050 187.345 ;
        RECT 76.140 186.905 78.050 187.205 ;
        RECT 76.140 186.090 76.440 186.905 ;
        RECT 77.460 186.695 78.050 186.905 ;
        RECT 95.750 186.090 96.050 188.880 ;
        RECT 76.140 185.790 96.050 186.090 ;
        RECT 76.140 185.785 76.440 185.790 ;
        RECT 96.650 185.110 96.950 191.695 ;
        RECT 98.735 191.555 99.325 191.695 ;
        RECT 104.360 189.715 104.960 211.245 ;
        RECT 105.230 212.955 107.605 213.095 ;
        RECT 105.230 205.900 105.370 212.955 ;
        RECT 107.015 212.700 107.605 212.955 ;
        RECT 113.740 211.770 114.440 213.765 ;
        RECT 112.445 211.070 114.440 211.770 ;
        RECT 105.565 210.220 106.165 210.860 ;
        RECT 106.720 206.910 107.310 207.560 ;
        RECT 107.015 205.900 107.605 206.155 ;
        RECT 105.230 205.760 107.605 205.900 ;
        RECT 105.230 198.995 105.370 205.760 ;
        RECT 107.015 205.505 107.605 205.760 ;
        RECT 113.740 205.005 114.440 211.070 ;
        RECT 112.445 204.305 114.440 205.005 ;
        RECT 105.565 203.140 106.165 203.780 ;
        RECT 106.805 199.845 107.395 200.495 ;
        RECT 107.015 198.995 107.605 199.250 ;
        RECT 105.230 198.855 107.605 198.995 ;
        RECT 105.230 192.015 105.370 198.855 ;
        RECT 107.015 198.600 107.605 198.855 ;
        RECT 112.390 197.810 113.090 197.870 ;
        RECT 113.740 197.810 114.440 204.305 ;
        RECT 112.390 197.110 114.440 197.810 ;
        RECT 105.565 196.270 106.165 196.910 ;
        RECT 106.805 192.965 107.395 193.615 ;
        RECT 107.015 192.015 107.605 192.270 ;
        RECT 105.230 191.875 107.605 192.015 ;
        RECT 97.370 188.930 97.970 189.570 ;
        RECT 102.885 185.805 103.475 186.455 ;
        RECT 105.230 185.110 105.370 191.875 ;
        RECT 107.015 191.620 107.605 191.875 ;
        RECT 113.740 190.390 114.440 197.110 ;
        RECT 119.930 190.390 124.435 214.945 ;
        RECT 112.445 189.690 124.435 190.390 ;
        RECT 105.565 188.930 106.165 189.570 ;
        RECT 106.805 185.805 107.395 186.455 ;
        RECT 96.650 184.810 119.510 185.110 ;
        RECT 56.400 183.815 64.115 184.115 ;
        RECT 56.400 183.650 56.980 183.815 ;
        RECT 58.295 181.180 58.525 183.040 ;
        RECT 118.630 182.840 118.860 183.040 ;
        RECT 119.210 182.840 119.510 184.810 ;
        RECT 118.630 182.700 119.510 182.840 ;
        RECT 118.630 182.390 118.860 182.700 ;
        RECT 58.295 178.760 58.525 180.620 ;
        RECT 118.630 179.970 118.860 181.830 ;
        RECT 58.295 176.340 58.525 178.200 ;
        RECT 118.630 177.550 118.860 179.410 ;
        RECT 119.930 176.990 124.435 189.690 ;
        RECT 118.630 176.340 124.435 176.990 ;
        RECT 54.935 174.845 88.470 175.545 ;
        RECT 53.610 173.975 54.200 174.625 ;
        RECT 52.600 172.655 53.190 172.835 ;
        RECT 53.755 172.655 54.055 173.975 ;
        RECT 52.600 172.355 54.055 172.655 ;
        RECT 52.600 172.185 53.190 172.355 ;
        RECT 37.435 171.070 46.490 171.115 ;
        RECT 37.435 170.420 46.915 171.070 ;
        RECT 37.435 170.415 46.490 170.420 ;
        RECT 37.435 166.635 43.110 170.415 ;
        RECT 44.330 169.400 45.030 170.415 ;
        RECT 53.755 168.915 54.055 172.355 ;
        RECT 87.770 171.690 88.470 174.845 ;
        RECT 104.660 173.345 113.515 174.045 ;
        RECT 89.000 172.685 89.590 173.335 ;
        RECT 87.645 170.680 88.595 171.690 ;
        RECT 104.660 171.420 105.360 173.345 ;
        RECT 106.835 173.175 107.425 173.345 ;
        RECT 90.940 170.720 105.360 171.420 ;
        RECT 112.815 172.085 113.515 173.345 ;
        RECT 119.930 172.085 124.435 176.340 ;
        RECT 112.815 171.385 124.435 172.085 ;
        RECT 53.585 168.265 54.175 168.915 ;
        RECT 37.435 165.935 46.970 166.635 ;
        RECT 52.365 166.585 52.955 167.235 ;
        RECT 37.435 161.980 43.110 165.935 ;
        RECT 44.410 164.785 45.110 165.935 ;
        RECT 53.755 164.605 54.055 168.265 ;
        RECT 53.615 163.955 54.205 164.605 ;
        RECT 46.270 161.980 46.970 162.045 ;
        RECT 37.435 161.280 46.970 161.980 ;
        RECT 52.300 161.950 52.890 162.600 ;
        RECT 37.435 136.020 43.110 161.280 ;
        RECT 44.330 160.295 45.030 161.280 ;
        RECT 53.755 160.005 54.055 163.955 ;
        RECT 87.770 161.730 88.470 170.680 ;
        RECT 89.025 168.715 89.615 169.365 ;
        RECT 89.015 162.625 89.605 163.275 ;
        RECT 87.735 160.720 88.685 161.730 ;
        RECT 92.050 161.500 92.750 170.720 ;
        RECT 105.535 169.865 106.135 170.505 ;
        RECT 107.055 167.910 107.645 168.000 ;
        RECT 104.935 167.610 107.645 167.910 ;
        RECT 93.740 163.090 94.330 163.305 ;
        RECT 104.935 163.090 105.235 167.610 ;
        RECT 107.055 167.350 107.645 167.610 ;
        RECT 106.780 166.600 107.480 166.655 ;
        RECT 106.780 165.900 113.505 166.600 ;
        RECT 112.805 165.530 113.505 165.900 ;
        RECT 119.930 165.530 124.435 171.385 ;
        RECT 112.805 164.855 124.435 165.530 ;
        RECT 112.860 164.830 124.435 164.855 ;
        RECT 93.740 162.790 105.235 163.090 ;
        RECT 105.535 163.075 106.135 163.715 ;
        RECT 93.740 162.655 94.330 162.790 ;
        RECT 90.950 160.800 92.750 161.500 ;
        RECT 104.935 160.695 105.235 162.790 ;
        RECT 107.055 160.695 107.645 160.870 ;
        RECT 104.935 160.395 107.645 160.695 ;
        RECT 107.055 160.220 107.645 160.395 ;
        RECT 53.595 159.355 54.185 160.005 ;
        RECT 85.885 159.215 86.500 159.220 ;
        RECT 85.850 157.850 86.500 159.215 ;
        RECT 89.025 158.725 89.615 159.375 ;
        RECT 52.305 157.200 52.895 157.850 ;
        RECT 55.245 157.150 113.390 157.850 ;
        RECT 85.850 157.140 86.500 157.150 ;
        RECT 112.690 155.380 113.390 157.150 ;
        RECT 45.655 153.520 45.885 155.380 ;
        RECT 110.660 154.730 113.390 155.380 ;
        RECT 45.655 151.100 45.885 152.960 ;
        RECT 110.660 152.310 110.890 154.170 ;
        RECT 45.655 148.680 45.885 150.540 ;
        RECT 110.660 149.890 110.890 151.750 ;
        RECT 45.655 146.260 45.885 148.120 ;
        RECT 110.660 147.470 110.890 149.330 ;
        RECT 45.655 143.840 45.885 145.700 ;
        RECT 110.660 145.050 110.890 146.910 ;
        RECT 45.655 141.420 45.885 143.280 ;
        RECT 110.660 142.630 110.890 144.490 ;
        RECT 112.690 142.955 113.390 154.730 ;
        RECT 45.655 139.000 45.885 140.860 ;
        RECT 110.660 140.210 110.890 142.070 ;
        RECT 45.655 136.580 45.885 138.440 ;
        RECT 110.660 137.790 110.890 139.650 ;
        RECT 110.660 136.580 111.960 137.230 ;
        RECT 111.310 136.020 111.960 136.580 ;
        RECT 37.435 135.370 111.960 136.020 ;
        RECT 37.435 135.055 43.110 135.370 ;
        RECT 112.435 135.055 117.435 142.955 ;
        RECT 119.930 135.055 124.435 164.830 ;
        RECT 114.575 122.715 115.575 135.055 ;
        RECT 30.605 110.755 36.715 111.565 ;
        RECT 10.695 109.755 36.715 110.755 ;
        RECT 125.980 110.355 130.860 111.565 ;
        RECT 30.605 89.350 36.715 109.755 ;
        RECT 45.870 109.315 46.770 109.475 ;
        RECT 54.855 109.325 55.755 109.485 ;
        RECT 65.090 109.325 65.990 109.485 ;
        RECT 45.850 108.675 46.790 109.315 ;
        RECT 54.835 108.685 55.775 109.325 ;
        RECT 65.070 108.685 66.010 109.325 ;
        RECT 73.495 109.300 74.075 109.940 ;
        RECT 78.595 109.850 79.495 110.010 ;
        RECT 45.870 108.515 46.770 108.675 ;
        RECT 54.855 108.525 55.755 108.685 ;
        RECT 65.090 108.525 65.990 108.685 ;
        RECT 44.115 106.800 45.015 106.960 ;
        RECT 44.095 106.160 45.035 106.800 ;
        RECT 61.330 106.655 62.230 106.815 ;
        RECT 71.355 106.655 72.255 106.815 ;
        RECT 44.115 106.000 45.015 106.160 ;
        RECT 51.565 105.865 52.155 106.515 ;
        RECT 61.310 106.015 62.250 106.655 ;
        RECT 71.335 106.015 72.275 106.655 ;
        RECT 73.605 106.310 73.745 109.300 ;
        RECT 78.575 109.210 79.515 109.850 ;
        RECT 125.980 109.355 134.175 110.355 ;
        RECT 78.595 109.050 79.495 109.210 ;
        RECT 81.780 107.735 82.360 107.920 ;
        RECT 125.980 107.735 130.860 109.355 ;
        RECT 81.735 107.035 130.860 107.735 ;
        RECT 45.795 102.330 46.795 103.330 ;
        RECT 45.870 100.465 46.770 100.625 ;
        RECT 45.850 99.825 46.790 100.465 ;
        RECT 45.870 99.665 46.770 99.825 ;
        RECT 51.805 97.640 51.945 105.865 ;
        RECT 61.330 105.855 62.230 106.015 ;
        RECT 71.355 105.855 72.255 106.015 ;
        RECT 73.365 105.660 73.955 106.310 ;
        RECT 82.185 106.030 82.765 106.225 ;
        RECT 82.185 105.890 83.135 106.030 ;
        RECT 54.005 103.900 54.595 104.550 ;
        RECT 51.790 97.440 51.945 97.640 ;
        RECT 44.115 97.005 45.015 97.165 ;
        RECT 44.095 96.365 45.035 97.005 ;
        RECT 51.790 96.405 51.930 97.440 ;
        RECT 44.115 96.205 45.015 96.365 ;
        RECT 51.585 95.755 52.175 96.405 ;
        RECT 45.795 92.420 46.795 93.420 ;
        RECT 37.195 89.350 37.775 89.600 ;
        RECT 30.605 89.210 37.775 89.350 ;
        RECT 45.870 89.245 46.770 89.405 ;
        RECT 30.605 58.355 36.715 89.210 ;
        RECT 37.195 88.960 37.775 89.210 ;
        RECT 45.850 88.605 46.790 89.245 ;
        RECT 45.870 88.445 46.770 88.605 ;
        RECT 44.115 87.645 45.015 87.805 ;
        RECT 44.095 87.005 45.035 87.645 ;
        RECT 44.115 86.845 45.015 87.005 ;
        RECT 51.790 86.330 51.930 95.755 ;
        RECT 54.230 94.620 54.370 103.900 ;
        RECT 64.165 103.870 64.755 104.520 ;
        RECT 54.780 102.365 55.780 103.365 ;
        RECT 64.385 100.190 64.525 103.870 ;
        RECT 65.275 102.305 66.275 103.305 ;
        RECT 73.605 102.975 73.745 105.660 ;
        RECT 82.185 105.585 82.765 105.890 ;
        RECT 82.995 105.085 83.135 105.890 ;
        RECT 82.940 104.435 83.170 105.085 ;
        RECT 74.215 102.975 75.165 103.345 ;
        RECT 73.605 102.835 75.165 102.975 ;
        RECT 79.245 102.940 80.145 103.100 ;
        RECT 73.605 100.190 73.745 102.835 ;
        RECT 74.215 102.335 75.165 102.835 ;
        RECT 79.225 102.300 80.165 102.940 ;
        RECT 79.245 102.140 80.145 102.300 ;
        RECT 82.940 102.015 83.170 103.875 ;
        RECT 123.775 103.225 124.005 105.085 ;
        RECT 64.385 100.050 73.745 100.190 ;
        RECT 54.855 99.365 55.755 99.525 ;
        RECT 54.835 98.725 55.775 99.365 ;
        RECT 54.855 98.565 55.755 98.725 ;
        RECT 64.385 98.325 64.525 100.050 ;
        RECT 65.090 99.385 65.990 99.545 ;
        RECT 65.070 98.745 66.010 99.385 ;
        RECT 65.090 98.585 65.990 98.745 ;
        RECT 64.165 97.675 64.755 98.325 ;
        RECT 61.330 96.305 62.230 96.465 ;
        RECT 61.310 95.665 62.250 96.305 ;
        RECT 61.330 95.505 62.230 95.665 ;
        RECT 54.005 93.970 54.595 94.620 ;
        RECT 51.565 85.680 52.155 86.330 ;
        RECT 45.795 82.265 46.795 83.265 ;
        RECT 45.870 80.170 46.770 80.330 ;
        RECT 45.850 79.530 46.790 80.170 ;
        RECT 45.870 79.370 46.770 79.530 ;
        RECT 43.510 77.160 44.410 77.320 ;
        RECT 43.490 76.520 44.430 77.160 ;
        RECT 51.790 77.130 51.930 85.680 ;
        RECT 54.230 84.570 54.370 93.970 ;
        RECT 54.780 92.455 55.780 93.455 ;
        RECT 54.855 89.595 55.755 89.755 ;
        RECT 54.835 88.955 55.775 89.595 ;
        RECT 54.855 88.795 55.755 88.955 ;
        RECT 64.385 88.320 64.525 97.675 ;
        RECT 71.355 96.305 72.255 96.465 ;
        RECT 73.605 96.345 73.745 100.050 ;
        RECT 78.520 99.850 79.420 100.010 ;
        RECT 78.500 99.210 79.440 99.850 ;
        RECT 82.940 99.595 83.170 101.455 ;
        RECT 123.775 100.805 124.005 102.665 ;
        RECT 125.980 100.250 130.860 107.035 ;
        RECT 123.900 100.245 130.860 100.250 ;
        RECT 123.775 99.595 130.860 100.245 ;
        RECT 123.900 99.550 130.860 99.595 ;
        RECT 78.520 99.050 79.420 99.210 ;
        RECT 125.980 99.050 130.860 99.550 ;
        RECT 122.020 98.350 130.860 99.050 ;
        RECT 93.345 97.875 112.655 98.015 ;
        RECT 71.335 95.665 72.275 96.305 ;
        RECT 73.385 95.695 73.975 96.345 ;
        RECT 93.345 96.285 93.485 97.875 ;
        RECT 112.515 96.880 112.655 97.875 ;
        RECT 93.230 96.015 93.820 96.285 ;
        RECT 86.065 95.875 93.820 96.015 ;
        RECT 71.355 95.505 72.255 95.665 ;
        RECT 65.275 92.410 66.275 93.410 ;
        RECT 73.605 92.965 73.745 95.695 ;
        RECT 74.215 92.965 75.165 93.445 ;
        RECT 79.245 93.420 80.145 93.580 ;
        RECT 73.605 92.825 75.165 92.965 ;
        RECT 65.090 89.720 65.990 89.880 ;
        RECT 65.070 89.080 66.010 89.720 ;
        RECT 65.090 88.920 65.990 89.080 ;
        RECT 64.165 87.670 64.755 88.320 ;
        RECT 61.330 86.285 62.230 86.445 ;
        RECT 61.310 85.645 62.250 86.285 ;
        RECT 61.330 85.485 62.230 85.645 ;
        RECT 54.005 83.920 54.595 84.570 ;
        RECT 54.220 80.980 54.360 83.920 ;
        RECT 54.780 82.440 55.780 83.440 ;
        RECT 64.390 80.980 64.530 87.670 ;
        RECT 71.355 86.445 72.255 86.605 ;
        RECT 73.605 86.585 73.745 92.825 ;
        RECT 74.215 92.435 75.165 92.825 ;
        RECT 79.225 92.780 80.165 93.420 ;
        RECT 79.245 92.620 80.145 92.780 ;
        RECT 78.520 90.020 79.420 90.180 ;
        RECT 78.500 89.380 79.440 90.020 ;
        RECT 78.520 89.220 79.420 89.380 ;
        RECT 71.335 85.805 72.275 86.445 ;
        RECT 73.325 85.935 73.915 86.585 ;
        RECT 71.355 85.645 72.255 85.805 ;
        RECT 73.605 84.680 73.745 85.935 ;
        RECT 73.590 84.540 73.745 84.680 ;
        RECT 65.275 82.555 66.275 83.555 ;
        RECT 54.220 80.840 64.530 80.980 ;
        RECT 54.220 79.150 54.360 80.840 ;
        RECT 54.855 80.160 55.755 80.320 ;
        RECT 54.835 79.520 55.775 80.160 ;
        RECT 54.855 79.360 55.755 79.520 ;
        RECT 54.005 78.500 54.595 79.150 ;
        RECT 64.390 79.055 64.530 80.840 ;
        RECT 65.090 80.205 65.990 80.365 ;
        RECT 65.070 79.565 66.010 80.205 ;
        RECT 65.090 79.405 65.990 79.565 ;
        RECT 64.165 78.405 64.755 79.055 ;
        RECT 61.330 77.350 62.230 77.510 ;
        RECT 51.585 76.865 52.175 77.130 ;
        RECT 52.360 76.865 52.940 77.115 ;
        RECT 51.585 76.725 52.940 76.865 ;
        RECT 43.510 76.360 44.410 76.520 ;
        RECT 51.585 76.480 52.175 76.725 ;
        RECT 52.360 76.475 52.940 76.725 ;
        RECT 61.310 76.710 62.250 77.350 ;
        RECT 71.355 77.120 72.255 77.280 ;
        RECT 61.330 76.550 62.230 76.710 ;
        RECT 71.335 76.480 72.275 77.120 ;
        RECT 73.605 76.885 73.745 84.540 ;
        RECT 74.320 82.705 75.320 83.705 ;
        RECT 79.210 83.065 80.110 83.225 ;
        RECT 79.190 82.425 80.130 83.065 ;
        RECT 79.210 82.265 80.110 82.425 ;
        RECT 78.680 79.895 79.580 80.055 ;
        RECT 78.660 79.255 79.600 79.895 ;
        RECT 78.680 79.095 79.580 79.255 ;
        RECT 86.065 77.270 86.205 95.875 ;
        RECT 93.230 95.635 93.820 95.875 ;
        RECT 96.465 95.630 97.465 96.630 ;
        RECT 97.970 96.255 98.870 96.415 ;
        RECT 97.950 95.615 98.890 96.255 ;
        RECT 112.265 96.230 112.855 96.880 ;
        RECT 114.795 95.630 115.795 96.630 ;
        RECT 116.300 96.255 117.200 96.415 ;
        RECT 116.280 95.615 117.220 96.255 ;
        RECT 97.970 95.455 98.870 95.615 ;
        RECT 116.300 95.455 117.200 95.615 ;
        RECT 96.040 95.005 96.940 95.165 ;
        RECT 114.370 95.005 115.270 95.165 ;
        RECT 94.560 93.905 95.560 94.905 ;
        RECT 96.020 94.365 96.960 95.005 ;
        RECT 96.040 94.205 96.940 94.365 ;
        RECT 93.530 92.340 94.530 93.340 ;
        RECT 94.990 93.335 95.890 93.495 ;
        RECT 94.970 92.695 95.910 93.335 ;
        RECT 104.595 93.220 105.595 94.220 ;
        RECT 112.890 93.905 113.890 94.905 ;
        RECT 114.350 94.365 115.290 95.005 ;
        RECT 114.370 94.205 115.270 94.365 ;
        RECT 94.990 92.535 95.890 92.695 ;
        RECT 111.860 92.340 112.860 93.340 ;
        RECT 113.320 93.335 114.220 93.495 ;
        RECT 113.300 92.695 114.240 93.335 ;
        RECT 113.320 92.535 114.220 92.695 ;
        RECT 89.675 90.940 90.575 91.100 ;
        RECT 89.655 90.300 90.595 90.940 ;
        RECT 91.180 90.835 92.180 91.835 ;
        RECT 92.875 91.755 93.775 91.915 ;
        RECT 92.855 91.115 93.795 91.755 ;
        RECT 92.875 90.955 93.775 91.115 ;
        RECT 108.005 90.940 108.905 91.100 ;
        RECT 107.985 90.300 108.925 90.940 ;
        RECT 109.510 90.835 110.510 91.835 ;
        RECT 111.205 91.755 112.105 91.915 ;
        RECT 111.185 91.115 112.125 91.755 ;
        RECT 111.205 90.955 112.105 91.115 ;
        RECT 89.675 90.140 90.575 90.300 ;
        RECT 108.005 90.140 108.905 90.300 ;
        RECT 87.965 88.675 88.965 89.675 ;
        RECT 89.675 88.580 90.575 88.740 ;
        RECT 106.295 88.695 107.295 89.695 ;
        RECT 125.980 89.650 130.860 98.350 ;
        RECT 121.885 88.950 130.860 89.650 ;
        RECT 108.005 88.580 108.905 88.740 ;
        RECT 89.655 87.940 90.595 88.580 ;
        RECT 107.985 87.940 108.925 88.580 ;
        RECT 89.675 87.780 90.575 87.940 ;
        RECT 108.005 87.780 108.905 87.940 ;
        RECT 90.500 86.295 91.500 87.295 ;
        RECT 92.010 87.115 92.910 87.275 ;
        RECT 91.990 86.475 92.930 87.115 ;
        RECT 92.010 86.315 92.910 86.475 ;
        RECT 108.830 86.295 109.830 87.295 ;
        RECT 110.340 87.115 111.240 87.275 ;
        RECT 110.320 86.475 111.260 87.115 ;
        RECT 110.340 86.315 111.240 86.475 ;
        RECT 92.575 84.870 93.575 85.870 ;
        RECT 94.115 85.595 95.015 85.755 ;
        RECT 94.095 84.955 95.035 85.595 ;
        RECT 94.115 84.795 95.015 84.955 ;
        RECT 110.905 84.870 111.905 85.870 ;
        RECT 112.445 85.595 113.345 85.755 ;
        RECT 112.425 84.955 113.365 85.595 ;
        RECT 112.445 84.795 113.345 84.955 ;
        RECT 92.575 82.925 93.575 83.925 ;
        RECT 94.320 83.770 95.220 83.930 ;
        RECT 94.300 83.130 95.240 83.770 ;
        RECT 94.320 82.970 95.220 83.130 ;
        RECT 110.905 82.925 111.905 83.925 ;
        RECT 112.650 83.770 113.550 83.930 ;
        RECT 112.630 83.130 113.570 83.770 ;
        RECT 112.650 82.970 113.550 83.130 ;
        RECT 94.845 81.385 95.845 82.385 ;
        RECT 96.400 82.310 97.300 82.470 ;
        RECT 96.380 81.670 97.320 82.310 ;
        RECT 96.400 81.510 97.300 81.670 ;
        RECT 98.000 81.385 99.000 82.385 ;
        RECT 113.175 81.385 114.175 82.385 ;
        RECT 114.730 82.310 115.630 82.470 ;
        RECT 114.710 81.670 115.650 82.310 ;
        RECT 114.730 81.510 115.630 81.670 ;
        RECT 116.330 81.385 117.330 82.385 ;
        RECT 93.095 79.035 111.935 79.175 ;
        RECT 93.095 77.900 93.235 79.035 ;
        RECT 92.920 77.270 93.510 77.900 ;
        RECT 96.225 77.340 97.225 78.340 ;
        RECT 97.680 77.965 98.580 78.125 ;
        RECT 97.660 77.325 98.600 77.965 ;
        RECT 111.795 77.525 111.935 79.035 ;
        RECT 86.065 77.250 93.510 77.270 ;
        RECT 86.065 77.130 93.235 77.250 ;
        RECT 97.680 77.165 98.580 77.325 ;
        RECT 71.355 76.320 72.255 76.480 ;
        RECT 73.345 76.235 73.935 76.885 ;
        RECT 45.795 73.260 46.795 74.260 ;
        RECT 54.780 73.235 55.780 74.235 ;
        RECT 65.275 73.380 66.275 74.380 ;
        RECT 73.915 73.080 74.915 74.080 ;
        RECT 79.340 73.545 80.240 73.705 ;
        RECT 79.320 72.905 80.260 73.545 ;
        RECT 79.340 72.745 80.240 72.905 ;
        RECT 51.555 72.165 52.455 72.325 ;
        RECT 51.535 71.525 52.475 72.165 ;
        RECT 51.555 71.365 52.455 71.525 ;
        RECT 58.280 69.580 58.860 70.220 ;
        RECT 58.465 68.875 58.605 69.580 ;
        RECT 74.370 69.410 74.950 69.660 ;
        RECT 75.630 69.410 76.220 69.665 ;
        RECT 63.550 69.195 64.450 69.355 ;
        RECT 74.370 69.270 76.220 69.410 ;
        RECT 58.240 68.225 58.830 68.875 ;
        RECT 63.530 68.555 64.470 69.195 ;
        RECT 74.370 69.020 74.950 69.270 ;
        RECT 75.630 69.015 76.220 69.270 ;
        RECT 63.550 68.395 64.450 68.555 ;
        RECT 51.390 66.060 52.390 67.060 ;
        RECT 51.555 65.625 52.455 65.785 ;
        RECT 51.535 64.985 52.475 65.625 ;
        RECT 51.555 64.825 52.455 64.985 ;
        RECT 58.480 63.540 58.620 68.225 ;
        RECT 63.550 67.375 64.450 67.535 ;
        RECT 63.530 66.735 64.470 67.375 ;
        RECT 75.855 67.150 75.995 69.015 ;
        RECT 63.550 66.575 64.450 66.735 ;
        RECT 75.630 66.500 76.220 67.150 ;
        RECT 63.550 65.555 64.450 65.715 ;
        RECT 63.530 64.915 64.470 65.555 ;
        RECT 63.550 64.755 64.450 64.915 ;
        RECT 75.855 64.545 75.995 66.500 ;
        RECT 63.560 63.740 64.460 63.900 ;
        RECT 75.630 63.895 76.220 64.545 ;
        RECT 58.260 62.890 58.850 63.540 ;
        RECT 63.540 63.100 64.480 63.740 ;
        RECT 63.560 62.940 64.460 63.100 ;
        RECT 47.840 59.955 48.420 60.185 ;
        RECT 45.150 59.815 48.420 59.955 ;
        RECT 30.605 58.340 37.710 58.355 ;
        RECT 30.605 57.700 38.000 58.340 ;
        RECT 30.605 57.655 37.710 57.700 ;
        RECT 30.605 47.680 36.715 57.655 ;
        RECT 30.605 46.980 38.000 47.680 ;
        RECT 30.605 46.125 36.715 46.980 ;
        RECT 37.230 46.125 38.540 46.470 ;
        RECT 30.605 45.425 38.540 46.125 ;
        RECT 43.645 45.700 44.545 45.860 ;
        RECT 30.605 39.545 36.715 45.425 ;
        RECT 37.230 45.100 38.540 45.425 ;
        RECT 43.625 45.060 44.565 45.700 ;
        RECT 43.645 44.900 44.545 45.060 ;
        RECT 45.150 43.325 45.290 59.815 ;
        RECT 47.840 59.545 48.420 59.815 ;
        RECT 51.390 59.370 52.390 60.370 ;
        RECT 51.555 58.930 52.455 59.090 ;
        RECT 51.535 58.290 52.475 58.930 ;
        RECT 51.555 58.130 52.455 58.290 ;
        RECT 58.465 55.055 58.605 62.890 ;
        RECT 63.560 61.915 64.460 62.075 ;
        RECT 75.855 62.015 75.995 63.895 ;
        RECT 63.540 61.275 64.480 61.915 ;
        RECT 75.630 61.365 76.220 62.015 ;
        RECT 63.560 61.115 64.460 61.275 ;
        RECT 63.560 60.090 64.460 60.250 ;
        RECT 63.540 59.450 64.480 60.090 ;
        RECT 63.560 59.290 64.460 59.450 ;
        RECT 75.855 59.370 75.995 61.365 ;
        RECT 75.630 58.720 76.220 59.370 ;
        RECT 63.550 58.280 64.450 58.440 ;
        RECT 63.530 57.640 64.470 58.280 ;
        RECT 63.550 57.480 64.450 57.640 ;
        RECT 75.855 56.895 75.995 58.720 ;
        RECT 61.255 56.455 62.155 56.615 ;
        RECT 63.560 56.455 64.460 56.615 ;
        RECT 61.235 55.815 62.175 56.455 ;
        RECT 63.540 55.815 64.480 56.455 ;
        RECT 75.630 56.245 76.220 56.895 ;
        RECT 73.050 55.970 73.630 56.235 ;
        RECT 74.305 55.970 74.895 56.225 ;
        RECT 73.050 55.830 74.895 55.970 ;
        RECT 61.255 55.655 62.155 55.815 ;
        RECT 63.560 55.655 64.460 55.815 ;
        RECT 73.050 55.595 73.630 55.830 ;
        RECT 74.305 55.575 74.895 55.830 ;
        RECT 86.065 55.500 86.205 77.130 ;
        RECT 111.570 76.875 112.160 77.525 ;
        RECT 114.825 77.095 115.825 78.095 ;
        RECT 116.330 77.720 117.230 77.880 ;
        RECT 116.310 77.080 117.250 77.720 ;
        RECT 116.330 76.920 117.230 77.080 ;
        RECT 95.750 76.715 96.650 76.875 ;
        RECT 94.270 75.615 95.270 76.615 ;
        RECT 95.730 76.075 96.670 76.715 ;
        RECT 114.400 76.470 115.300 76.630 ;
        RECT 95.750 75.915 96.650 76.075 ;
        RECT 112.920 75.370 113.920 76.370 ;
        RECT 114.380 75.830 115.320 76.470 ;
        RECT 114.400 75.670 115.300 75.830 ;
        RECT 93.240 74.050 94.240 75.050 ;
        RECT 94.700 75.045 95.600 75.205 ;
        RECT 94.680 74.405 95.620 75.045 ;
        RECT 94.700 74.245 95.600 74.405 ;
        RECT 111.890 73.805 112.890 74.805 ;
        RECT 113.350 74.800 114.250 74.960 ;
        RECT 113.330 74.160 114.270 74.800 ;
        RECT 113.350 74.000 114.250 74.160 ;
        RECT 89.385 72.650 90.285 72.810 ;
        RECT 89.365 72.010 90.305 72.650 ;
        RECT 90.890 72.545 91.890 73.545 ;
        RECT 92.585 73.465 93.485 73.625 ;
        RECT 92.565 72.825 93.505 73.465 ;
        RECT 92.585 72.665 93.485 72.825 ;
        RECT 108.035 72.405 108.935 72.565 ;
        RECT 89.385 71.850 90.285 72.010 ;
        RECT 108.015 71.765 108.955 72.405 ;
        RECT 109.540 72.300 110.540 73.300 ;
        RECT 111.235 73.220 112.135 73.380 ;
        RECT 111.215 72.580 112.155 73.220 ;
        RECT 111.235 72.420 112.135 72.580 ;
        RECT 108.035 71.605 108.935 71.765 ;
        RECT 87.675 70.405 88.675 71.405 ;
        RECT 89.385 70.290 90.285 70.450 ;
        RECT 89.365 69.650 90.305 70.290 ;
        RECT 106.325 70.175 107.325 71.175 ;
        RECT 125.980 71.045 130.860 88.950 ;
        RECT 122.170 70.345 130.860 71.045 ;
        RECT 108.035 70.045 108.935 70.205 ;
        RECT 89.385 69.490 90.285 69.650 ;
        RECT 108.015 69.405 108.955 70.045 ;
        RECT 108.035 69.245 108.935 69.405 ;
        RECT 90.210 68.005 91.210 69.005 ;
        RECT 91.720 68.825 92.620 68.985 ;
        RECT 91.700 68.185 92.640 68.825 ;
        RECT 91.720 68.025 92.620 68.185 ;
        RECT 108.860 67.760 109.860 68.760 ;
        RECT 110.370 68.580 111.270 68.740 ;
        RECT 110.350 67.940 111.290 68.580 ;
        RECT 110.370 67.780 111.270 67.940 ;
        RECT 92.285 66.580 93.285 67.580 ;
        RECT 93.825 67.305 94.725 67.465 ;
        RECT 93.805 66.665 94.745 67.305 ;
        RECT 93.825 66.505 94.725 66.665 ;
        RECT 110.935 66.335 111.935 67.335 ;
        RECT 112.475 67.060 113.375 67.220 ;
        RECT 112.455 66.420 113.395 67.060 ;
        RECT 112.475 66.260 113.375 66.420 ;
        RECT 92.285 64.635 93.285 65.635 ;
        RECT 94.030 65.480 94.930 65.640 ;
        RECT 94.010 64.840 94.950 65.480 ;
        RECT 104.070 65.290 104.660 65.665 ;
        RECT 94.030 64.680 94.930 64.840 ;
        RECT 94.555 63.095 95.555 64.095 ;
        RECT 96.110 64.020 97.010 64.180 ;
        RECT 96.090 63.380 97.030 64.020 ;
        RECT 96.110 63.220 97.010 63.380 ;
        RECT 97.710 63.095 98.710 64.095 ;
        RECT 104.015 61.200 104.715 65.290 ;
        RECT 110.935 64.390 111.935 65.390 ;
        RECT 112.680 65.235 113.580 65.395 ;
        RECT 112.660 64.595 113.600 65.235 ;
        RECT 112.680 64.435 113.580 64.595 ;
        RECT 113.205 62.850 114.205 63.850 ;
        RECT 114.760 63.775 115.660 63.935 ;
        RECT 114.740 63.135 115.680 63.775 ;
        RECT 114.760 62.975 115.660 63.135 ;
        RECT 116.360 62.850 117.360 63.850 ;
        RECT 125.980 61.200 130.860 70.345 ;
        RECT 104.015 60.500 130.860 61.200 ;
        RECT 104.045 59.830 104.745 60.500 ;
        RECT 75.765 55.360 86.205 55.500 ;
        RECT 101.560 59.130 104.745 59.830 ;
        RECT 58.240 54.405 58.830 55.055 ;
        RECT 75.765 55.020 75.905 55.360 ;
        RECT 60.340 54.880 75.905 55.020 ;
        RECT 51.390 52.705 52.390 53.705 ;
        RECT 51.480 52.000 52.380 52.160 ;
        RECT 51.460 51.360 52.400 52.000 ;
        RECT 51.480 51.200 52.380 51.360 ;
        RECT 58.480 49.485 58.620 54.405 ;
        RECT 60.340 52.870 60.480 54.880 ;
        RECT 101.560 54.235 102.260 59.130 ;
        RECT 107.025 58.145 107.925 58.305 ;
        RECT 107.005 57.505 107.945 58.145 ;
        RECT 107.025 57.345 107.925 57.505 ;
        RECT 108.560 57.215 109.560 58.215 ;
        RECT 110.030 58.145 110.930 58.305 ;
        RECT 110.010 57.505 110.950 58.145 ;
        RECT 110.030 57.345 110.930 57.505 ;
        RECT 111.560 57.215 112.560 58.215 ;
        RECT 114.000 58.145 114.900 58.305 ;
        RECT 113.980 57.505 114.920 58.145 ;
        RECT 114.000 57.345 114.900 57.505 ;
        RECT 106.310 55.805 107.310 56.805 ;
        RECT 71.810 53.535 102.260 54.235 ;
        RECT 105.975 54.130 106.975 55.130 ;
        RECT 107.580 55.070 108.480 55.230 ;
        RECT 107.560 54.430 108.500 55.070 ;
        RECT 107.580 54.270 108.480 54.430 ;
        RECT 59.990 51.860 60.940 52.870 ;
        RECT 63.785 52.490 64.685 52.650 ;
        RECT 60.395 50.310 60.535 51.860 ;
        RECT 63.765 51.850 64.705 52.490 ;
        RECT 73.050 52.190 73.630 52.485 ;
        RECT 74.670 52.190 75.260 52.445 ;
        RECT 73.050 52.050 75.260 52.190 ;
        RECT 61.405 50.815 62.405 51.815 ;
        RECT 63.785 51.690 64.685 51.850 ;
        RECT 73.050 51.845 73.630 52.050 ;
        RECT 74.670 51.795 75.260 52.050 ;
        RECT 75.575 52.045 76.275 53.535 ;
        RECT 106.540 52.895 107.440 53.055 ;
        RECT 106.520 52.255 107.460 52.895 ;
        RECT 106.540 52.095 107.440 52.255 ;
        RECT 75.515 51.765 76.275 52.045 ;
        RECT 75.515 51.625 76.390 51.765 ;
        RECT 125.980 51.755 130.860 60.500 ;
        RECT 75.515 51.345 76.275 51.625 ;
        RECT 63.785 50.670 64.685 50.830 ;
        RECT 60.100 49.670 60.680 50.310 ;
        RECT 63.765 50.030 64.705 50.670 ;
        RECT 58.260 48.835 58.850 49.485 ;
        RECT 61.405 48.930 62.405 49.930 ;
        RECT 63.785 49.870 64.685 50.030 ;
        RECT 72.940 49.930 73.940 50.930 ;
        RECT 75.780 49.455 75.920 51.345 ;
        RECT 105.975 50.510 106.975 51.510 ;
        RECT 121.810 51.055 130.860 51.755 ;
        RECT 106.540 49.615 107.440 49.775 ;
        RECT 63.785 48.850 64.685 49.010 ;
        RECT 63.765 48.210 64.705 48.850 ;
        RECT 75.555 48.805 76.145 49.455 ;
        RECT 106.520 48.975 107.460 49.615 ;
        RECT 106.540 48.815 107.440 48.975 ;
        RECT 61.405 47.105 62.405 48.105 ;
        RECT 63.785 48.050 64.685 48.210 ;
        RECT 72.880 47.360 73.880 48.360 ;
        RECT 51.390 46.080 52.390 47.080 ;
        RECT 63.795 47.030 64.695 47.190 ;
        RECT 63.775 46.390 64.715 47.030 ;
        RECT 75.775 46.900 75.915 48.805 ;
        RECT 63.795 46.230 64.695 46.390 ;
        RECT 75.550 46.250 76.140 46.900 ;
        RECT 105.975 46.760 106.975 47.760 ;
        RECT 107.580 47.575 108.480 47.735 ;
        RECT 107.560 46.935 108.500 47.575 ;
        RECT 107.580 46.775 108.480 46.935 ;
        RECT 48.220 45.695 49.120 45.855 ;
        RECT 48.200 45.055 49.140 45.695 ;
        RECT 61.405 45.230 62.405 46.230 ;
        RECT 63.795 45.210 64.695 45.370 ;
        RECT 48.220 44.895 49.120 45.055 ;
        RECT 63.775 44.570 64.715 45.210 ;
        RECT 72.990 44.855 73.990 45.855 ;
        RECT 63.795 44.410 64.695 44.570 ;
        RECT 46.720 43.555 47.620 43.715 ;
        RECT 44.960 42.675 45.550 43.325 ;
        RECT 46.700 42.915 47.640 43.555 ;
        RECT 61.405 43.410 62.405 44.410 ;
        RECT 75.815 44.335 75.955 46.250 ;
        RECT 106.650 45.155 107.650 46.155 ;
        RECT 107.580 44.445 108.480 44.605 ;
        RECT 75.590 43.685 76.180 44.335 ;
        RECT 107.560 43.805 108.500 44.445 ;
        RECT 63.795 43.385 64.695 43.545 ;
        RECT 46.720 42.755 47.620 42.915 ;
        RECT 39.315 39.850 40.315 40.850 ;
        RECT 37.230 39.545 38.540 39.740 ;
        RECT 30.605 38.845 38.540 39.545 ;
        RECT 43.665 39.040 44.565 39.200 ;
        RECT 30.605 33.050 36.715 38.845 ;
        RECT 37.230 38.370 38.540 38.845 ;
        RECT 43.645 38.400 44.585 39.040 ;
        RECT 43.665 38.240 44.565 38.400 ;
        RECT 45.150 37.250 45.290 42.675 ;
        RECT 55.020 42.260 55.610 42.910 ;
        RECT 63.775 42.745 64.715 43.385 ;
        RECT 48.125 39.860 49.125 40.860 ;
        RECT 48.220 39.065 49.120 39.225 ;
        RECT 48.200 38.425 49.140 39.065 ;
        RECT 48.220 38.265 49.120 38.425 ;
        RECT 55.260 37.250 55.400 42.260 ;
        RECT 61.405 41.670 62.405 42.670 ;
        RECT 63.795 42.585 64.695 42.745 ;
        RECT 72.990 42.245 73.990 43.245 ;
        RECT 75.790 41.775 75.930 43.685 ;
        RECT 107.580 43.645 108.480 43.805 ;
        RECT 109.060 43.665 110.060 44.665 ;
        RECT 110.480 44.420 111.380 44.580 ;
        RECT 110.460 43.780 111.400 44.420 ;
        RECT 110.480 43.620 111.380 43.780 ;
        RECT 111.790 43.705 112.790 44.705 ;
        RECT 114.000 44.675 114.900 44.835 ;
        RECT 113.980 44.035 114.920 44.675 ;
        RECT 125.980 44.655 130.860 51.055 ;
        RECT 125.705 44.605 130.860 44.655 ;
        RECT 114.000 43.875 114.900 44.035 ;
        RECT 125.340 43.965 130.860 44.605 ;
        RECT 125.705 43.955 130.860 43.965 ;
        RECT 63.785 41.575 64.685 41.735 ;
        RECT 63.765 40.935 64.705 41.575 ;
        RECT 75.565 41.125 76.155 41.775 ;
        RECT 97.185 41.145 98.185 42.145 ;
        RECT 112.745 41.615 113.335 42.265 ;
        RECT 61.405 39.835 62.405 40.835 ;
        RECT 63.785 40.775 64.685 40.935 ;
        RECT 63.795 39.750 64.695 39.910 ;
        RECT 72.990 39.760 73.990 40.760 ;
        RECT 63.775 39.110 64.715 39.750 ;
        RECT 63.795 38.950 64.695 39.110 ;
        RECT 73.085 38.725 73.665 38.895 ;
        RECT 70.055 38.425 74.680 38.725 ;
        RECT 45.150 37.105 45.295 37.250 ;
        RECT 55.260 37.105 55.405 37.250 ;
        RECT 45.155 36.620 45.295 37.105 ;
        RECT 44.930 35.970 45.520 36.620 ;
        RECT 46.720 36.590 47.620 36.750 ;
        RECT 37.230 33.050 38.540 33.645 ;
        RECT 38.965 33.145 39.965 34.145 ;
        RECT 30.605 32.350 38.540 33.050 ;
        RECT 43.625 32.925 44.525 33.085 ;
        RECT 30.605 26.825 36.715 32.350 ;
        RECT 37.230 32.275 38.540 32.350 ;
        RECT 43.605 32.285 44.545 32.925 ;
        RECT 43.625 32.125 44.525 32.285 ;
        RECT 45.155 30.530 45.295 35.970 ;
        RECT 46.700 35.950 47.640 36.590 ;
        RECT 55.265 36.575 55.405 37.105 ;
        RECT 57.680 37.000 58.580 37.160 ;
        RECT 46.720 35.790 47.620 35.950 ;
        RECT 55.040 35.925 55.630 36.575 ;
        RECT 57.660 36.360 58.600 37.000 ;
        RECT 57.680 36.200 58.580 36.360 ;
        RECT 48.110 33.155 49.110 34.155 ;
        RECT 49.410 32.905 50.310 33.065 ;
        RECT 49.390 32.265 50.330 32.905 ;
        RECT 49.410 32.105 50.310 32.265 ;
        RECT 55.265 30.550 55.405 35.925 ;
        RECT 58.965 35.625 59.965 36.625 ;
        RECT 66.580 34.865 67.170 34.925 ;
        RECT 66.580 34.275 67.310 34.865 ;
        RECT 58.965 32.580 59.965 33.580 ;
        RECT 44.930 29.880 45.520 30.530 ;
        RECT 46.720 30.305 47.620 30.465 ;
        RECT 37.400 26.825 38.710 27.275 ;
        RECT 38.965 27.030 39.965 28.030 ;
        RECT 30.605 26.125 38.710 26.825 ;
        RECT 43.665 26.500 44.565 26.660 ;
        RECT 30.605 18.240 36.715 26.125 ;
        RECT 37.400 25.905 38.710 26.125 ;
        RECT 43.645 25.860 44.585 26.500 ;
        RECT 43.665 25.700 44.565 25.860 ;
        RECT 45.155 24.055 45.295 29.880 ;
        RECT 46.700 29.665 47.640 30.305 ;
        RECT 55.040 29.900 55.630 30.550 ;
        RECT 46.720 29.505 47.620 29.665 ;
        RECT 48.145 27.060 49.145 28.060 ;
        RECT 49.410 26.500 50.310 26.660 ;
        RECT 49.390 25.860 50.330 26.500 ;
        RECT 49.410 25.700 50.310 25.860 ;
        RECT 46.720 24.230 47.620 24.390 ;
        RECT 44.930 23.405 45.520 24.055 ;
        RECT 46.700 23.590 47.640 24.230 ;
        RECT 55.265 24.205 55.405 29.900 ;
        RECT 56.890 27.590 63.725 28.240 ;
        RECT 46.720 23.430 47.620 23.590 ;
        RECT 55.040 23.555 55.630 24.205 ;
        RECT 37.975 20.635 38.975 21.635 ;
        RECT 45.155 19.170 45.295 23.405 ;
        RECT 48.100 20.655 49.100 21.655 ;
        RECT 55.265 19.170 55.405 23.555 ;
        RECT 45.155 19.030 55.405 19.170 ;
        RECT 56.890 18.240 57.540 27.590 ;
        RECT 63.495 25.170 63.725 27.030 ;
        RECT 63.495 22.750 63.725 24.610 ;
        RECT 30.605 17.590 57.540 18.240 ;
        RECT 30.605 11.775 36.715 17.590 ;
        RECT 66.610 17.040 67.310 34.275 ;
        RECT 70.055 33.375 70.355 38.425 ;
        RECT 73.085 38.255 73.665 38.425 ;
        RECT 74.380 37.515 74.680 38.425 ;
        RECT 75.735 38.095 75.875 41.125 ;
        RECT 76.040 38.095 76.630 38.350 ;
        RECT 75.735 37.955 76.630 38.095 ;
        RECT 76.040 37.700 76.630 37.955 ;
        RECT 72.830 35.980 73.780 36.990 ;
        RECT 74.315 36.875 74.895 37.515 ;
        RECT 70.760 35.085 71.660 35.245 ;
        RECT 70.740 34.445 71.680 35.085 ;
        RECT 70.760 34.285 71.660 34.445 ;
        RECT 73.295 33.375 73.885 33.560 ;
        RECT 70.055 33.075 73.885 33.375 ;
        RECT 73.295 32.910 73.885 33.075 ;
        RECT 57.335 11.760 67.335 17.040 ;
        RECT 80.565 16.855 81.265 35.115 ;
        RECT 88.560 26.380 88.790 28.240 ;
        RECT 88.560 23.960 88.790 25.820 ;
        RECT 88.560 22.750 89.770 23.400 ;
        RECT 89.120 19.610 89.770 22.750 ;
        RECT 97.335 19.785 98.035 41.145 ;
        RECT 112.970 40.785 113.110 41.615 ;
        RECT 112.670 40.145 113.250 40.785 ;
        RECT 97.185 19.610 98.185 19.785 ;
        RECT 89.120 18.960 98.185 19.610 ;
        RECT 89.120 17.025 89.770 18.960 ;
        RECT 97.185 18.785 98.185 18.960 ;
        RECT 71.275 11.780 81.275 16.855 ;
        RECT 88.240 11.785 98.240 17.025 ;
        RECT 65.365 6.335 66.365 11.760 ;
        RECT 79.725 8.425 80.725 11.780 ;
        RECT 96.915 10.700 97.915 11.785 ;
        RECT 125.980 11.775 130.860 43.955 ;
        RECT 96.915 9.700 155.690 10.700 ;
        RECT 154.575 8.955 155.690 9.700 ;
        RECT 154.575 8.905 155.670 8.955 ;
        RECT 79.725 7.425 135.355 8.425 ;
        RECT 65.365 5.335 113.245 6.335 ;
      LAYER met2 ;
        RECT 56.935 219.630 58.105 219.645 ;
        RECT 56.925 218.630 60.880 219.630 ;
        RECT 56.935 218.515 58.105 218.630 ;
        RECT 132.095 215.945 133.265 215.990 ;
        RECT 127.560 214.945 133.265 215.945 ;
        RECT 132.095 214.860 133.265 214.945 ;
        RECT 7.795 214.715 8.965 214.730 ;
        RECT 7.785 213.715 11.740 214.715 ;
        RECT 7.795 213.600 8.965 213.715 ;
        RECT 97.305 210.015 98.035 210.785 ;
        RECT 105.500 210.155 106.230 210.925 ;
        RECT 102.805 207.455 103.385 207.555 ;
        RECT 106.725 207.455 107.305 207.555 ;
        RECT 63.855 207.175 64.435 207.345 ;
        RECT 92.940 207.175 93.520 207.345 ;
        RECT 102.805 207.315 107.305 207.455 ;
        RECT 63.855 206.875 95.050 207.175 ;
        RECT 102.805 206.915 103.385 207.315 ;
        RECT 63.855 206.705 64.435 206.875 ;
        RECT 92.940 206.705 93.520 206.875 ;
        RECT 53.280 206.215 53.860 206.415 ;
        RECT 53.280 205.915 60.585 206.215 ;
        RECT 53.280 205.775 53.860 205.915 ;
        RECT 53.240 201.375 53.820 201.605 ;
        RECT 60.285 201.375 60.585 205.915 ;
        RECT 63.675 203.390 64.255 203.540 ;
        RECT 92.940 203.390 93.520 203.560 ;
        RECT 63.675 203.090 93.520 203.390 ;
        RECT 63.675 202.900 64.255 203.090 ;
        RECT 92.940 202.920 93.520 203.090 ;
        RECT 63.815 202.425 64.115 202.900 ;
        RECT 63.675 201.785 64.255 202.425 ;
        RECT 53.240 201.075 76.390 201.375 ;
        RECT 53.240 200.965 53.820 201.075 ;
        RECT 76.090 198.135 76.390 201.075 ;
        RECT 75.990 197.495 76.570 198.135 ;
        RECT 52.950 186.535 54.080 187.705 ;
        RECT 56.400 183.650 56.980 184.290 ;
        RECT 54.215 181.770 54.795 181.940 ;
        RECT 56.545 181.770 56.845 183.650 ;
        RECT 54.215 181.470 56.845 181.770 ;
        RECT 54.215 181.300 54.795 181.470 ;
        RECT 89.005 173.160 89.585 173.330 ;
        RECT 89.005 173.120 93.305 173.160 ;
        RECT 94.750 173.120 95.050 206.875 ;
        RECT 97.305 202.840 98.035 203.610 ;
        RECT 102.890 200.240 103.470 200.490 ;
        RECT 105.035 200.240 105.175 207.315 ;
        RECT 106.725 206.915 107.305 207.315 ;
        RECT 105.500 203.075 106.230 203.845 ;
        RECT 106.810 200.240 107.390 200.490 ;
        RECT 102.890 200.100 107.390 200.240 ;
        RECT 102.890 199.850 103.470 200.100 ;
        RECT 97.305 195.890 98.035 196.660 ;
        RECT 102.890 193.360 103.470 193.610 ;
        RECT 105.035 193.360 105.175 200.100 ;
        RECT 106.810 199.850 107.390 200.100 ;
        RECT 105.500 196.205 106.230 196.975 ;
        RECT 106.810 193.360 107.390 193.610 ;
        RECT 102.890 193.220 107.390 193.360 ;
        RECT 102.890 192.970 103.470 193.220 ;
        RECT 95.535 188.815 96.265 189.585 ;
        RECT 97.305 188.865 98.035 189.635 ;
        RECT 97.305 186.200 98.035 186.605 ;
        RECT 102.890 186.200 103.470 186.450 ;
        RECT 105.035 186.200 105.175 193.220 ;
        RECT 106.810 192.970 107.390 193.220 ;
        RECT 105.500 188.865 106.230 189.635 ;
        RECT 106.810 186.200 107.390 186.450 ;
        RECT 97.305 186.060 107.390 186.200 ;
        RECT 97.305 185.835 98.035 186.060 ;
        RECT 102.890 185.810 103.470 186.060 ;
        RECT 106.810 185.810 107.390 186.060 ;
        RECT 89.005 172.860 95.050 173.120 ;
        RECT 89.005 172.690 89.585 172.860 ;
        RECT 93.005 172.820 95.050 172.860 ;
        RECT 89.030 169.145 89.610 169.360 ;
        RECT 85.990 168.845 89.610 169.145 ;
        RECT 52.515 167.270 53.215 167.275 ;
        RECT 52.285 166.570 55.005 167.270 ;
        RECT 52.305 162.590 52.885 162.595 ;
        RECT 54.305 162.590 55.005 166.570 ;
        RECT 52.305 161.955 55.005 162.590 ;
        RECT 52.345 161.890 55.005 161.955 ;
        RECT 52.310 157.830 53.205 157.845 ;
        RECT 54.305 157.830 55.005 161.890 ;
        RECT 85.990 159.215 86.290 168.845 ;
        RECT 89.030 168.720 89.610 168.845 ;
        RECT 89.020 163.100 89.600 163.270 ;
        RECT 93.005 163.100 93.305 172.820 ;
        RECT 105.470 169.800 106.200 170.570 ;
        RECT 93.745 163.100 94.325 163.300 ;
        RECT 89.020 162.800 94.325 163.100 ;
        RECT 105.470 163.010 106.200 163.780 ;
        RECT 89.020 162.630 89.600 162.800 ;
        RECT 93.745 162.660 94.325 162.800 ;
        RECT 85.885 159.200 86.465 159.215 ;
        RECT 89.030 159.200 89.610 159.370 ;
        RECT 85.885 158.900 89.610 159.200 ;
        RECT 85.885 158.575 86.465 158.900 ;
        RECT 89.030 158.730 89.610 158.900 ;
        RECT 55.185 157.830 55.885 157.845 ;
        RECT 52.250 157.130 55.885 157.830 ;
        RECT 111.295 123.665 112.465 123.725 ;
        RECT 111.295 122.665 115.555 123.665 ;
        RECT 111.295 122.595 112.465 122.665 ;
        RECT 7.795 110.805 8.965 110.820 ;
        RECT 7.785 109.805 11.740 110.805 ;
        RECT 137.750 110.355 138.920 110.400 ;
        RECT 53.975 110.200 82.835 110.340 ;
        RECT 7.795 109.690 8.965 109.805 ;
        RECT 45.870 109.285 46.770 109.475 ;
        RECT 43.415 108.585 46.770 109.285 ;
        RECT 43.415 106.960 44.115 108.585 ;
        RECT 45.870 108.515 46.770 108.585 ;
        RECT 53.975 109.075 54.115 110.200 ;
        RECT 54.855 109.075 55.755 109.485 ;
        RECT 53.975 108.935 55.755 109.075 ;
        RECT 43.415 106.000 45.015 106.960 ;
        RECT 43.415 100.610 44.115 106.000 ;
        RECT 45.730 102.245 46.860 103.415 ;
        RECT 45.870 100.610 46.770 100.625 ;
        RECT 43.415 99.910 46.770 100.610 ;
        RECT 43.415 97.165 44.115 99.910 ;
        RECT 45.740 99.875 46.770 99.910 ;
        RECT 45.870 99.665 46.770 99.875 ;
        RECT 53.975 99.025 54.115 108.935 ;
        RECT 54.855 108.525 55.755 108.935 ;
        RECT 64.160 109.075 64.300 110.200 ;
        RECT 65.090 109.075 65.990 109.485 ;
        RECT 73.420 109.235 74.150 110.005 ;
        RECT 78.595 109.950 79.495 110.010 ;
        RECT 78.595 109.250 81.550 109.950 ;
        RECT 64.160 108.935 65.990 109.075 ;
        RECT 78.595 109.050 79.495 109.250 ;
        RECT 61.330 106.685 62.230 106.815 ;
        RECT 61.310 105.855 62.230 106.685 ;
        RECT 54.715 102.280 55.845 103.450 ;
        RECT 54.855 99.025 55.755 99.525 ;
        RECT 53.965 98.885 55.755 99.025 ;
        RECT 43.415 96.205 45.015 97.165 ;
        RECT 37.195 89.590 37.775 89.600 ;
        RECT 43.415 89.590 44.115 96.205 ;
        RECT 45.730 92.335 46.860 93.505 ;
        RECT 37.195 89.405 46.320 89.590 ;
        RECT 37.195 88.960 46.770 89.405 ;
        RECT 53.975 89.345 54.115 98.885 ;
        RECT 54.855 98.565 55.755 98.885 ;
        RECT 61.310 96.465 62.010 105.855 ;
        RECT 64.160 99.045 64.300 108.935 ;
        RECT 65.090 108.525 65.990 108.935 ;
        RECT 80.850 107.995 81.550 109.250 ;
        RECT 80.850 107.295 82.420 107.995 ;
        RECT 71.355 105.855 72.255 106.815 ;
        RECT 65.210 102.220 66.340 103.390 ;
        RECT 65.090 99.045 65.990 99.545 ;
        RECT 64.160 98.905 65.990 99.045 ;
        RECT 61.310 95.505 62.230 96.465 ;
        RECT 54.715 92.370 55.845 93.540 ;
        RECT 54.855 89.345 55.755 89.755 ;
        RECT 53.965 89.205 55.755 89.345 ;
        RECT 37.485 88.890 46.770 88.960 ;
        RECT 43.415 87.805 44.115 88.890 ;
        RECT 45.870 88.445 46.770 88.890 ;
        RECT 43.415 86.845 45.015 87.805 ;
        RECT 43.415 80.160 44.115 86.845 ;
        RECT 45.730 82.180 46.860 83.350 ;
        RECT 45.870 80.160 46.770 80.330 ;
        RECT 43.415 79.460 46.770 80.160 ;
        RECT 53.975 79.880 54.115 89.205 ;
        RECT 54.855 88.795 55.755 89.205 ;
        RECT 61.310 86.445 62.010 95.505 ;
        RECT 64.160 89.470 64.300 98.905 ;
        RECT 65.090 98.585 65.990 98.905 ;
        RECT 71.455 96.465 72.155 105.855 ;
        RECT 79.245 102.970 80.145 103.100 ;
        RECT 79.230 102.140 80.145 102.970 ;
        RECT 79.230 102.000 79.930 102.140 ;
        RECT 80.850 102.000 81.550 107.295 ;
        RECT 81.720 107.280 82.420 107.295 ;
        RECT 82.695 106.225 82.835 110.200 ;
        RECT 133.215 109.355 138.920 110.355 ;
        RECT 137.750 109.270 138.920 109.355 ;
        RECT 82.185 105.835 82.835 106.225 ;
        RECT 82.185 105.585 82.765 105.835 ;
        RECT 78.590 101.300 81.550 102.000 ;
        RECT 78.590 100.010 79.290 101.300 ;
        RECT 78.520 99.050 79.420 100.010 ;
        RECT 71.355 95.505 72.255 96.465 ;
        RECT 65.210 92.325 66.340 93.495 ;
        RECT 65.090 89.470 65.990 89.880 ;
        RECT 64.160 89.330 65.990 89.470 ;
        RECT 61.310 85.485 62.230 86.445 ;
        RECT 54.715 82.355 55.845 83.525 ;
        RECT 54.855 79.880 55.755 80.320 ;
        RECT 53.975 79.740 55.755 79.880 ;
        RECT 43.415 77.320 44.115 79.460 ;
        RECT 45.870 79.370 46.770 79.460 ;
        RECT 54.855 79.360 55.755 79.740 ;
        RECT 61.310 77.510 62.010 85.485 ;
        RECT 64.160 79.910 64.300 89.330 ;
        RECT 65.090 88.920 65.990 89.330 ;
        RECT 71.455 86.605 72.155 95.505 ;
        RECT 79.245 92.620 80.145 93.580 ;
        RECT 79.345 91.725 80.045 92.620 ;
        RECT 80.850 91.725 81.550 101.300 ;
        RECT 121.955 98.315 122.685 99.085 ;
        RECT 95.945 97.175 116.800 97.315 ;
        RECT 95.945 95.165 96.085 97.175 ;
        RECT 96.400 95.545 97.530 96.715 ;
        RECT 98.290 96.415 98.430 97.175 ;
        RECT 97.970 95.455 98.870 96.415 ;
        RECT 94.495 93.820 95.625 94.990 ;
        RECT 95.945 94.615 96.940 95.165 ;
        RECT 96.040 94.205 96.940 94.615 ;
        RECT 78.565 91.025 81.550 91.725 ;
        RECT 90.055 92.600 92.970 92.740 ;
        RECT 90.055 91.100 90.195 92.600 ;
        RECT 78.565 90.180 79.265 91.025 ;
        RECT 78.520 89.220 79.420 90.180 ;
        RECT 71.355 85.645 72.255 86.605 ;
        RECT 65.210 82.470 66.340 83.640 ;
        RECT 65.090 79.910 65.990 80.365 ;
        RECT 64.160 79.770 65.990 79.910 ;
        RECT 65.090 79.405 65.990 79.770 ;
        RECT 43.415 76.490 44.410 77.320 ;
        RECT 43.510 76.360 44.410 76.490 ;
        RECT 52.285 76.410 53.015 77.180 ;
        RECT 61.310 76.550 62.230 77.510 ;
        RECT 71.455 77.280 72.155 85.645 ;
        RECT 74.255 82.620 75.385 83.790 ;
        RECT 79.210 82.265 80.110 83.225 ;
        RECT 79.385 81.530 80.085 82.265 ;
        RECT 80.850 81.530 81.550 91.025 ;
        RECT 89.675 90.140 90.575 91.100 ;
        RECT 91.115 90.750 92.245 91.920 ;
        RECT 92.830 91.915 92.970 92.600 ;
        RECT 93.465 92.255 94.595 93.425 ;
        RECT 94.990 93.085 95.890 93.495 ;
        RECT 96.330 93.085 96.470 94.205 ;
        RECT 94.990 92.945 96.470 93.085 ;
        RECT 94.990 92.535 95.890 92.945 ;
        RECT 92.830 91.700 93.775 91.915 ;
        RECT 95.370 91.700 95.510 92.535 ;
        RECT 92.830 91.560 95.510 91.700 ;
        RECT 92.830 91.365 93.775 91.560 ;
        RECT 92.875 90.955 93.775 91.365 ;
        RECT 87.900 88.590 89.030 89.760 ;
        RECT 90.055 88.740 90.195 90.140 ;
        RECT 89.675 88.330 90.575 88.740 ;
        RECT 89.635 87.780 90.575 88.330 ;
        RECT 89.635 85.550 89.775 87.780 ;
        RECT 90.435 86.210 91.565 87.380 ;
        RECT 92.010 86.830 92.910 87.275 ;
        RECT 92.010 86.690 94.635 86.830 ;
        RECT 92.010 86.315 92.910 86.690 ;
        RECT 92.155 85.550 92.295 86.315 ;
        RECT 89.635 85.410 92.295 85.550 ;
        RECT 91.650 82.270 91.790 85.410 ;
        RECT 92.510 84.785 93.640 85.955 ;
        RECT 94.495 85.755 94.635 86.690 ;
        RECT 94.115 84.795 95.015 85.755 ;
        RECT 92.510 82.840 93.640 84.010 ;
        RECT 94.320 83.520 95.220 83.930 ;
        RECT 94.235 82.970 95.220 83.520 ;
        RECT 94.235 82.270 94.375 82.970 ;
        RECT 91.650 82.130 94.375 82.270 ;
        RECT 78.750 80.830 81.550 81.530 ;
        RECT 78.750 80.055 79.450 80.830 ;
        RECT 78.680 79.095 79.580 80.055 ;
        RECT 45.730 73.175 46.860 74.345 ;
        RECT 54.715 73.150 55.845 74.320 ;
        RECT 51.555 72.305 52.455 72.325 ;
        RECT 50.825 72.165 52.455 72.305 ;
        RECT 50.825 65.740 50.965 72.165 ;
        RECT 51.555 71.365 52.455 72.165 ;
        RECT 61.310 71.315 62.010 76.550 ;
        RECT 71.355 76.320 72.255 77.280 ;
        RECT 65.210 73.295 66.340 74.465 ;
        RECT 71.455 71.315 72.155 76.320 ;
        RECT 73.850 72.995 74.980 74.165 ;
        RECT 79.340 72.745 80.240 73.705 ;
        RECT 79.505 71.315 80.205 72.745 ;
        RECT 80.850 71.315 81.550 80.830 ;
        RECT 93.300 80.530 93.440 82.130 ;
        RECT 94.780 81.300 95.910 82.470 ;
        RECT 96.400 81.510 97.300 82.470 ;
        RECT 96.780 80.530 96.920 81.510 ;
        RECT 97.935 81.300 99.065 82.470 ;
        RECT 93.300 80.390 96.920 80.530 ;
        RECT 104.045 78.780 104.185 97.175 ;
        RECT 114.275 95.165 114.415 97.175 ;
        RECT 114.730 95.545 115.860 96.715 ;
        RECT 116.660 96.415 116.800 97.175 ;
        RECT 116.300 95.455 117.200 96.415 ;
        RECT 104.530 93.135 105.660 94.305 ;
        RECT 112.825 93.820 113.955 94.990 ;
        RECT 114.275 94.615 115.270 95.165 ;
        RECT 114.370 94.205 115.270 94.615 ;
        RECT 108.385 92.600 111.300 92.740 ;
        RECT 108.385 91.100 108.525 92.600 ;
        RECT 108.005 90.140 108.905 91.100 ;
        RECT 109.445 90.750 110.575 91.920 ;
        RECT 111.160 91.915 111.300 92.600 ;
        RECT 111.795 92.255 112.925 93.425 ;
        RECT 113.320 93.085 114.220 93.495 ;
        RECT 114.660 93.085 114.800 94.205 ;
        RECT 113.320 92.945 114.800 93.085 ;
        RECT 113.320 92.535 114.220 92.945 ;
        RECT 111.160 91.700 112.105 91.915 ;
        RECT 113.700 91.700 113.840 92.535 ;
        RECT 111.160 91.560 113.840 91.700 ;
        RECT 111.160 91.365 112.105 91.560 ;
        RECT 111.205 90.955 112.105 91.365 ;
        RECT 106.230 88.610 107.360 89.780 ;
        RECT 108.385 88.740 108.525 90.140 ;
        RECT 108.005 88.330 108.905 88.740 ;
        RECT 107.965 87.780 108.905 88.330 ;
        RECT 107.965 85.550 108.105 87.780 ;
        RECT 108.765 86.210 109.895 87.380 ;
        RECT 110.340 86.830 111.240 87.275 ;
        RECT 110.340 86.690 112.965 86.830 ;
        RECT 110.340 86.315 111.240 86.690 ;
        RECT 110.485 85.550 110.625 86.315 ;
        RECT 107.965 85.410 110.625 85.550 ;
        RECT 109.980 82.270 110.120 85.410 ;
        RECT 110.840 84.785 111.970 85.955 ;
        RECT 112.825 85.755 112.965 86.690 ;
        RECT 112.445 84.795 113.345 85.755 ;
        RECT 110.840 82.840 111.970 84.010 ;
        RECT 112.650 83.520 113.550 83.930 ;
        RECT 112.565 82.970 113.550 83.520 ;
        RECT 112.565 82.270 112.705 82.970 ;
        RECT 109.980 82.130 112.705 82.270 ;
        RECT 111.630 80.530 111.770 82.130 ;
        RECT 113.110 81.300 114.240 82.470 ;
        RECT 114.730 81.510 115.630 82.470 ;
        RECT 115.110 80.530 115.250 81.510 ;
        RECT 116.265 81.300 117.395 82.470 ;
        RECT 111.630 80.390 115.250 80.530 ;
        RECT 95.870 78.640 116.790 78.780 ;
        RECT 95.870 76.875 96.010 78.640 ;
        RECT 96.160 77.255 97.290 78.425 ;
        RECT 97.885 78.125 98.025 78.640 ;
        RECT 97.680 77.165 98.580 78.125 ;
        RECT 94.205 75.530 95.335 76.700 ;
        RECT 95.750 75.915 96.650 76.875 ;
        RECT 114.305 76.630 114.445 78.640 ;
        RECT 114.760 77.010 115.890 78.180 ;
        RECT 116.650 77.880 116.790 78.640 ;
        RECT 116.330 76.920 117.230 77.880 ;
        RECT 89.765 74.310 92.680 74.450 ;
        RECT 89.765 72.810 89.905 74.310 ;
        RECT 89.385 71.850 90.285 72.810 ;
        RECT 90.825 72.460 91.955 73.630 ;
        RECT 92.540 73.625 92.680 74.310 ;
        RECT 93.175 73.965 94.305 75.135 ;
        RECT 94.700 74.795 95.600 75.205 ;
        RECT 96.040 74.795 96.180 75.915 ;
        RECT 112.855 75.285 113.985 76.455 ;
        RECT 114.305 76.080 115.300 76.630 ;
        RECT 114.400 75.670 115.300 76.080 ;
        RECT 94.700 74.655 96.180 74.795 ;
        RECT 94.700 74.245 95.600 74.655 ;
        RECT 92.540 73.410 93.485 73.625 ;
        RECT 95.080 73.410 95.220 74.245 ;
        RECT 92.540 73.270 95.220 73.410 ;
        RECT 108.415 74.065 111.330 74.205 ;
        RECT 92.540 73.075 93.485 73.270 ;
        RECT 92.585 72.665 93.485 73.075 ;
        RECT 108.415 72.565 108.555 74.065 ;
        RECT 61.310 70.615 81.550 71.315 ;
        RECT 58.205 69.515 58.935 70.285 ;
        RECT 62.935 68.945 63.075 70.615 ;
        RECT 63.550 68.945 64.450 69.355 ;
        RECT 74.310 69.020 75.010 70.615 ;
        RECT 87.610 70.320 88.740 71.490 ;
        RECT 89.765 70.450 89.905 71.850 ;
        RECT 108.035 71.605 108.935 72.565 ;
        RECT 109.475 72.215 110.605 73.385 ;
        RECT 111.190 73.380 111.330 74.065 ;
        RECT 111.825 73.720 112.955 74.890 ;
        RECT 113.350 74.550 114.250 74.960 ;
        RECT 114.690 74.550 114.830 75.670 ;
        RECT 113.350 74.410 114.830 74.550 ;
        RECT 113.350 74.000 114.250 74.410 ;
        RECT 111.190 73.165 112.135 73.380 ;
        RECT 113.730 73.165 113.870 74.000 ;
        RECT 111.190 73.025 113.870 73.165 ;
        RECT 111.190 72.830 112.135 73.025 ;
        RECT 111.235 72.420 112.135 72.830 ;
        RECT 89.385 70.040 90.285 70.450 ;
        RECT 106.260 70.090 107.390 71.260 ;
        RECT 108.415 70.205 108.555 71.605 ;
        RECT 89.345 69.490 90.285 70.040 ;
        RECT 108.035 69.795 108.935 70.205 ;
        RECT 62.935 68.805 64.450 68.945 ;
        RECT 51.325 65.975 52.455 67.145 ;
        RECT 62.935 66.975 63.075 68.805 ;
        RECT 63.550 68.395 64.450 68.805 ;
        RECT 63.550 66.975 64.450 67.535 ;
        RECT 62.935 66.835 64.450 66.975 ;
        RECT 89.345 66.885 89.485 69.490 ;
        RECT 107.995 69.245 108.935 69.795 ;
        RECT 90.145 67.920 91.275 69.090 ;
        RECT 91.720 68.165 92.620 68.985 ;
        RECT 91.720 68.025 94.345 68.165 ;
        RECT 91.865 66.885 92.005 68.025 ;
        RECT 51.555 65.740 52.455 65.785 ;
        RECT 50.825 65.600 52.455 65.740 ;
        RECT 47.765 59.480 48.495 60.250 ;
        RECT 50.825 59.020 50.965 65.600 ;
        RECT 51.555 64.825 52.455 65.600 ;
        RECT 62.935 65.325 63.075 66.835 ;
        RECT 63.550 66.575 64.450 66.835 ;
        RECT 85.270 66.745 92.005 66.885 ;
        RECT 63.550 65.325 64.450 65.715 ;
        RECT 62.935 65.185 64.450 65.325 ;
        RECT 62.935 63.460 63.075 65.185 ;
        RECT 63.550 64.755 64.450 65.185 ;
        RECT 63.560 63.460 64.460 63.900 ;
        RECT 62.935 63.320 64.460 63.460 ;
        RECT 62.935 61.655 63.075 63.320 ;
        RECT 63.560 62.940 64.460 63.320 ;
        RECT 63.560 61.655 64.460 62.075 ;
        RECT 62.935 61.515 64.460 61.655 ;
        RECT 51.325 59.285 52.455 60.455 ;
        RECT 62.935 59.830 63.075 61.515 ;
        RECT 63.560 61.115 64.460 61.515 ;
        RECT 63.560 59.830 64.460 60.250 ;
        RECT 62.935 59.690 64.460 59.830 ;
        RECT 51.555 59.020 52.455 59.090 ;
        RECT 50.825 58.880 52.455 59.020 ;
        RECT 50.825 58.370 50.965 58.880 ;
        RECT 37.420 57.670 50.965 58.370 ;
        RECT 51.555 58.130 52.455 58.880 ;
        RECT 50.825 52.130 50.965 57.670 ;
        RECT 62.935 57.905 63.075 59.690 ;
        RECT 63.560 59.290 64.460 59.690 ;
        RECT 63.550 57.905 64.450 58.440 ;
        RECT 62.935 57.765 64.450 57.905 ;
        RECT 61.255 55.655 62.155 56.615 ;
        RECT 62.935 56.280 63.075 57.765 ;
        RECT 63.550 57.480 64.450 57.765 ;
        RECT 63.560 56.280 64.460 56.615 ;
        RECT 62.935 56.140 64.460 56.280 ;
        RECT 63.560 55.655 64.460 56.140 ;
        RECT 61.635 54.145 61.775 55.655 ;
        RECT 72.975 55.530 73.705 56.300 ;
        RECT 61.635 54.005 64.285 54.145 ;
        RECT 51.325 52.620 52.455 53.790 ;
        RECT 64.145 52.650 64.285 54.005 ;
        RECT 63.785 52.250 64.685 52.650 ;
        RECT 51.480 52.130 52.380 52.160 ;
        RECT 50.825 51.990 52.380 52.130 ;
        RECT 51.480 51.200 52.380 51.990 ;
        RECT 63.170 52.110 64.685 52.250 ;
        RECT 61.340 50.730 62.470 51.900 ;
        RECT 59.825 49.405 60.955 50.575 ;
        RECT 63.170 50.270 63.310 52.110 ;
        RECT 63.785 51.690 64.685 52.110 ;
        RECT 72.975 51.780 73.705 52.550 ;
        RECT 63.785 50.270 64.685 50.830 ;
        RECT 63.170 50.130 64.685 50.270 ;
        RECT 61.340 48.845 62.470 50.015 ;
        RECT 63.170 48.620 63.310 50.130 ;
        RECT 63.785 49.870 64.685 50.130 ;
        RECT 72.875 49.845 74.005 51.015 ;
        RECT 63.785 48.620 64.685 49.010 ;
        RECT 63.170 48.480 64.685 48.620 ;
        RECT 37.360 47.600 38.060 47.650 ;
        RECT 37.360 46.900 44.445 47.600 ;
        RECT 43.745 45.860 44.445 46.900 ;
        RECT 51.325 45.995 52.455 47.165 ;
        RECT 61.340 47.020 62.470 48.190 ;
        RECT 63.170 46.755 63.310 48.480 ;
        RECT 63.785 48.050 64.685 48.480 ;
        RECT 72.815 47.275 73.945 48.445 ;
        RECT 63.795 46.755 64.695 47.190 ;
        RECT 63.170 46.615 64.695 46.755 ;
        RECT 43.645 45.725 44.545 45.860 ;
        RECT 48.220 45.740 49.120 45.855 ;
        RECT 48.220 45.725 56.675 45.740 ;
        RECT 43.645 45.040 56.675 45.725 ;
        RECT 61.340 45.145 62.470 46.315 ;
        RECT 43.645 45.025 49.120 45.040 ;
        RECT 43.645 44.900 44.545 45.025 ;
        RECT 39.250 39.765 40.380 40.935 ;
        RECT 43.665 38.870 44.565 39.200 ;
        RECT 44.775 38.870 44.915 45.025 ;
        RECT 43.665 38.570 44.915 38.870 ;
        RECT 43.665 38.240 44.565 38.570 ;
        RECT 38.900 33.060 40.030 34.230 ;
        RECT 43.625 32.550 44.525 33.085 ;
        RECT 44.775 32.550 44.915 38.570 ;
        RECT 43.625 32.250 44.915 32.550 ;
        RECT 43.625 32.125 44.525 32.250 ;
        RECT 38.900 26.945 40.030 28.115 ;
        RECT 43.665 26.060 44.565 26.660 ;
        RECT 44.775 26.060 44.915 32.250 ;
        RECT 43.665 25.920 44.915 26.060 ;
        RECT 46.220 43.385 46.520 45.025 ;
        RECT 48.220 44.895 49.120 45.025 ;
        RECT 46.720 43.385 47.620 43.715 ;
        RECT 46.220 43.085 47.620 43.385 ;
        RECT 46.220 38.895 46.520 43.085 ;
        RECT 46.720 42.755 47.620 43.085 ;
        RECT 48.060 39.775 49.190 40.945 ;
        RECT 48.220 38.895 49.120 39.225 ;
        RECT 46.220 38.595 49.120 38.895 ;
        RECT 46.220 36.420 46.520 38.595 ;
        RECT 48.220 38.265 49.120 38.595 ;
        RECT 55.975 37.030 56.675 45.040 ;
        RECT 63.170 44.950 63.310 46.615 ;
        RECT 63.795 46.230 64.695 46.615 ;
        RECT 63.795 44.950 64.695 45.370 ;
        RECT 63.170 44.810 64.695 44.950 ;
        RECT 61.340 43.325 62.470 44.495 ;
        RECT 63.170 43.125 63.310 44.810 ;
        RECT 63.795 44.410 64.695 44.810 ;
        RECT 72.925 44.770 74.055 45.940 ;
        RECT 63.795 43.125 64.695 43.545 ;
        RECT 63.170 42.985 64.695 43.125 ;
        RECT 61.340 41.585 62.470 42.755 ;
        RECT 63.170 41.320 63.310 42.985 ;
        RECT 63.795 42.585 64.695 42.985 ;
        RECT 72.925 42.160 74.055 43.330 ;
        RECT 63.785 41.320 64.685 41.735 ;
        RECT 63.170 41.180 64.685 41.320 ;
        RECT 61.340 39.750 62.470 40.920 ;
        RECT 63.170 39.500 63.310 41.180 ;
        RECT 63.785 40.775 64.685 41.180 ;
        RECT 63.795 39.500 64.695 39.910 ;
        RECT 72.925 39.675 74.055 40.845 ;
        RECT 63.170 39.360 64.695 39.500 ;
        RECT 63.795 38.950 64.695 39.360 ;
        RECT 73.010 38.190 73.740 38.960 ;
        RECT 85.270 38.440 85.410 66.745 ;
        RECT 91.530 64.030 91.670 66.745 ;
        RECT 92.220 66.495 93.350 67.665 ;
        RECT 94.205 67.465 94.345 68.025 ;
        RECT 93.825 66.505 94.725 67.465 ;
        RECT 107.995 67.015 108.135 69.245 ;
        RECT 108.795 67.675 109.925 68.845 ;
        RECT 110.370 68.295 111.270 68.740 ;
        RECT 110.370 68.155 112.995 68.295 ;
        RECT 110.370 67.780 111.270 68.155 ;
        RECT 110.515 67.015 110.655 67.780 ;
        RECT 107.995 66.875 110.655 67.015 ;
        RECT 92.220 64.550 93.350 65.720 ;
        RECT 94.030 65.230 94.930 65.640 ;
        RECT 93.740 65.090 94.930 65.230 ;
        RECT 93.740 64.030 93.880 65.090 ;
        RECT 94.030 64.680 94.930 65.090 ;
        RECT 91.530 63.890 93.880 64.030 ;
        RECT 93.010 61.865 93.150 63.890 ;
        RECT 94.490 63.010 95.620 64.180 ;
        RECT 96.110 63.220 97.010 64.180 ;
        RECT 96.490 61.865 96.630 63.220 ;
        RECT 97.645 63.010 98.775 64.180 ;
        RECT 110.010 63.735 110.150 66.875 ;
        RECT 110.870 66.250 112.000 67.420 ;
        RECT 112.855 67.220 112.995 68.155 ;
        RECT 112.475 66.260 113.375 67.220 ;
        RECT 110.870 64.305 112.000 65.475 ;
        RECT 112.680 64.985 113.580 65.395 ;
        RECT 112.595 64.435 113.580 64.985 ;
        RECT 112.595 63.735 112.735 64.435 ;
        RECT 110.010 63.595 112.735 63.735 ;
        RECT 93.010 61.725 96.630 61.865 ;
        RECT 111.660 61.995 111.800 63.595 ;
        RECT 113.140 62.765 114.270 63.935 ;
        RECT 114.760 62.975 115.660 63.935 ;
        RECT 115.140 61.995 115.280 62.975 ;
        RECT 116.295 62.765 117.425 63.935 ;
        RECT 111.660 61.855 115.280 61.995 ;
        RECT 96.490 61.630 96.630 61.725 ;
        RECT 96.490 61.490 96.670 61.630 ;
        RECT 96.530 60.575 96.670 61.490 ;
        RECT 96.530 60.435 103.610 60.575 ;
        RECT 97.120 41.060 98.250 42.230 ;
        RECT 103.470 40.535 103.610 60.435 ;
        RECT 107.125 58.835 114.800 59.535 ;
        RECT 107.125 58.305 107.825 58.835 ;
        RECT 110.155 58.305 110.855 58.835 ;
        RECT 114.100 58.305 114.800 58.835 ;
        RECT 107.025 58.175 107.925 58.305 ;
        RECT 104.595 57.475 107.925 58.175 ;
        RECT 104.595 52.925 105.295 57.475 ;
        RECT 107.025 57.345 107.925 57.475 ;
        RECT 108.495 57.130 109.625 58.300 ;
        RECT 110.030 57.345 110.930 58.305 ;
        RECT 111.495 57.130 112.625 58.300 ;
        RECT 114.000 57.345 114.900 58.305 ;
        RECT 106.245 55.720 107.375 56.890 ;
        RECT 105.910 54.045 107.040 55.215 ;
        RECT 107.580 54.270 108.480 55.230 ;
        RECT 107.780 53.250 108.480 54.270 ;
        RECT 106.640 53.055 108.480 53.250 ;
        RECT 106.540 52.925 108.480 53.055 ;
        RECT 104.535 52.550 108.480 52.925 ;
        RECT 104.535 52.225 107.440 52.550 ;
        RECT 104.535 49.645 105.235 52.225 ;
        RECT 106.540 52.095 107.440 52.225 ;
        RECT 105.910 50.425 107.040 51.595 ;
        RECT 106.540 49.645 107.440 49.775 ;
        RECT 104.535 49.440 107.440 49.645 ;
        RECT 104.520 48.945 107.440 49.440 ;
        RECT 104.520 48.740 105.235 48.945 ;
        RECT 106.540 48.815 107.440 48.945 ;
        RECT 104.520 43.115 105.220 48.740 ;
        RECT 105.910 46.675 107.040 47.845 ;
        RECT 107.580 46.775 108.480 47.735 ;
        RECT 106.585 45.070 107.715 46.240 ;
        RECT 107.960 44.605 108.100 46.775 ;
        RECT 107.580 43.645 108.480 44.605 ;
        RECT 107.945 43.115 108.085 43.645 ;
        RECT 108.995 43.580 110.125 44.750 ;
        RECT 110.480 43.620 111.380 44.580 ;
        RECT 111.725 43.620 112.855 44.790 ;
        RECT 114.000 44.655 114.900 44.835 ;
        RECT 114.000 44.605 125.705 44.655 ;
        RECT 114.000 43.965 125.930 44.605 ;
        RECT 114.000 43.955 125.705 43.965 ;
        RECT 114.000 43.875 114.900 43.955 ;
        RECT 104.520 42.870 108.435 43.115 ;
        RECT 110.545 42.870 111.245 43.620 ;
        RECT 114.100 42.870 114.800 43.875 ;
        RECT 104.520 42.415 114.800 42.870 ;
        RECT 108.015 42.170 114.800 42.415 ;
        RECT 112.660 40.535 113.260 40.785 ;
        RECT 103.470 40.395 113.260 40.535 ;
        RECT 112.660 40.145 113.260 40.395 ;
        RECT 85.250 38.300 85.410 38.440 ;
        RECT 57.995 37.440 71.560 38.140 ;
        RECT 57.995 37.160 58.695 37.440 ;
        RECT 57.680 37.030 58.695 37.160 ;
        RECT 46.720 36.420 47.620 36.750 ;
        RECT 46.220 36.120 47.620 36.420 ;
        RECT 55.975 36.330 58.695 37.030 ;
        RECT 57.680 36.200 58.580 36.330 ;
        RECT 46.220 32.375 46.520 36.120 ;
        RECT 46.720 35.790 47.620 36.120 ;
        RECT 58.900 35.540 60.030 36.710 ;
        RECT 70.860 35.245 71.560 37.440 ;
        RECT 74.315 37.320 74.895 37.515 ;
        RECT 85.250 37.320 85.390 38.300 ;
        RECT 74.315 37.180 85.390 37.320 ;
        RECT 72.740 35.900 73.870 37.070 ;
        RECT 74.315 36.875 74.895 37.180 ;
        RECT 70.760 34.285 71.660 35.245 ;
        RECT 48.045 33.070 49.175 34.240 ;
        RECT 49.410 32.375 50.310 33.065 ;
        RECT 58.900 32.495 60.030 33.665 ;
        RECT 46.220 32.235 50.310 32.375 ;
        RECT 46.220 30.135 46.520 32.235 ;
        RECT 49.410 32.105 50.310 32.235 ;
        RECT 46.720 30.135 47.620 30.465 ;
        RECT 46.220 29.835 47.620 30.135 ;
        RECT 46.220 26.265 46.520 29.835 ;
        RECT 46.720 29.505 47.620 29.835 ;
        RECT 48.080 26.975 49.210 28.145 ;
        RECT 49.410 26.265 50.310 26.660 ;
        RECT 46.220 25.965 50.310 26.265 ;
        RECT 43.665 25.700 44.565 25.920 ;
        RECT 47.020 24.390 47.320 25.965 ;
        RECT 49.410 25.700 50.310 25.965 ;
        RECT 46.720 23.430 47.620 24.390 ;
        RECT 37.910 20.550 39.040 21.720 ;
        RECT 48.035 20.570 49.165 21.740 ;
        RECT 97.120 18.700 98.250 19.870 ;
        RECT 112.265 4.220 113.265 6.285 ;
        RECT 134.375 4.560 135.375 8.375 ;
        RECT 112.225 3.090 113.395 4.220 ;
        RECT 134.200 4.035 135.375 4.560 ;
        RECT 154.690 4.560 155.690 9.855 ;
        RECT 134.200 3.430 135.370 4.035 ;
        RECT 154.690 3.865 155.925 4.560 ;
        RECT 154.755 3.430 155.925 3.865 ;
      LAYER met3 ;
        RECT 56.935 219.640 58.105 219.645 ;
        RECT 56.930 218.520 58.110 219.640 ;
        RECT 56.935 218.515 58.105 218.520 ;
        RECT 132.095 215.985 133.265 215.990 ;
        RECT 132.090 214.865 133.270 215.985 ;
        RECT 132.095 214.860 133.265 214.865 ;
        RECT 7.795 214.725 8.965 214.730 ;
        RECT 7.790 213.605 8.970 214.725 ;
        RECT 7.795 213.600 8.965 213.605 ;
        RECT 97.520 210.785 97.820 210.790 ;
        RECT 97.305 210.015 98.035 210.785 ;
        RECT 105.500 210.155 106.230 210.925 ;
        RECT 97.520 206.615 97.820 210.015 ;
        RECT 105.715 206.615 106.015 210.155 ;
        RECT 97.520 206.315 106.015 206.615 ;
        RECT 97.520 203.610 97.820 206.315 ;
        RECT 105.715 203.845 106.015 206.315 ;
        RECT 97.305 202.840 98.035 203.610 ;
        RECT 105.500 203.075 106.230 203.845 ;
        RECT 97.520 196.660 97.820 202.840 ;
        RECT 105.715 196.975 106.015 203.075 ;
        RECT 97.305 195.890 98.035 196.660 ;
        RECT 105.500 196.205 106.230 196.975 ;
        RECT 97.520 189.635 97.820 195.890 ;
        RECT 105.715 189.635 106.015 196.205 ;
        RECT 95.535 189.350 96.265 189.585 ;
        RECT 97.305 189.350 98.035 189.635 ;
        RECT 95.535 189.050 98.035 189.350 ;
        RECT 95.535 188.815 96.265 189.050 ;
        RECT 97.305 188.865 98.035 189.050 ;
        RECT 105.500 188.865 106.230 189.635 ;
        RECT 52.950 187.205 54.080 187.705 ;
        RECT 52.950 186.905 57.225 187.205 ;
        RECT 52.950 186.535 54.080 186.905 ;
        RECT 56.925 185.405 57.225 186.905 ;
        RECT 97.305 185.835 98.035 186.605 ;
        RECT 97.520 185.405 97.820 185.835 ;
        RECT 56.925 185.105 97.820 185.405 ;
        RECT 105.715 170.570 106.015 188.865 ;
        RECT 105.470 169.800 106.200 170.570 ;
        RECT 105.715 163.780 106.015 169.800 ;
        RECT 105.470 163.010 106.200 163.780 ;
        RECT 111.295 123.720 112.465 123.725 ;
        RECT 111.290 122.600 112.470 123.720 ;
        RECT 111.295 122.595 112.465 122.600 ;
        RECT 7.795 110.815 8.965 110.820 ;
        RECT 7.790 109.695 8.970 110.815 ;
        RECT 137.750 110.395 138.920 110.400 ;
        RECT 73.420 109.885 74.150 110.005 ;
        RECT 44.060 109.870 74.150 109.885 ;
        RECT 7.795 109.690 8.965 109.695 ;
        RECT 42.710 109.585 74.150 109.870 ;
        RECT 42.710 109.570 44.360 109.585 ;
        RECT 42.710 102.665 43.010 109.570 ;
        RECT 73.420 109.235 74.150 109.585 ;
        RECT 137.745 109.275 138.925 110.395 ;
        RECT 137.750 109.270 138.920 109.275 ;
        RECT 45.730 102.665 46.860 103.415 ;
        RECT 42.710 102.365 46.860 102.665 ;
        RECT 42.710 92.795 43.010 102.365 ;
        RECT 45.730 102.245 46.860 102.365 ;
        RECT 54.715 102.280 55.845 103.450 ;
        RECT 55.130 100.775 55.430 102.280 ;
        RECT 65.210 102.220 66.340 103.390 ;
        RECT 65.395 101.200 65.695 102.220 ;
        RECT 53.465 100.475 55.430 100.775 ;
        RECT 63.830 100.900 65.775 101.200 ;
        RECT 45.730 92.795 46.860 93.505 ;
        RECT 42.710 92.495 46.860 92.795 ;
        RECT 45.730 92.335 46.860 92.495 ;
        RECT 53.465 93.215 53.765 100.475 ;
        RECT 54.715 93.215 55.845 93.540 ;
        RECT 53.465 92.915 55.845 93.215 ;
        RECT 45.730 82.700 46.860 83.350 ;
        RECT 44.765 82.400 46.860 82.700 ;
        RECT 44.765 73.790 45.065 82.400 ;
        RECT 45.730 82.180 46.860 82.400 ;
        RECT 53.465 83.090 53.765 92.915 ;
        RECT 54.715 92.370 55.845 92.915 ;
        RECT 63.830 92.935 64.130 100.900 ;
        RECT 121.955 99.050 122.685 99.085 ;
        RECT 104.705 98.350 122.685 99.050 ;
        RECT 96.400 96.520 97.530 96.715 ;
        RECT 94.710 95.820 97.530 96.520 ;
        RECT 94.710 94.990 95.410 95.820 ;
        RECT 96.400 95.545 97.530 95.820 ;
        RECT 94.495 94.765 95.625 94.990 ;
        RECT 93.375 94.065 95.625 94.765 ;
        RECT 104.705 94.305 105.405 98.350 ;
        RECT 121.955 98.315 122.685 98.350 ;
        RECT 114.730 96.520 115.860 96.715 ;
        RECT 113.040 95.820 115.860 96.520 ;
        RECT 113.040 94.990 113.740 95.820 ;
        RECT 114.730 95.545 115.860 95.820 ;
        RECT 112.825 94.765 113.955 94.990 ;
        RECT 65.210 92.935 66.340 93.495 ;
        RECT 93.375 93.425 94.075 94.065 ;
        RECT 94.495 93.820 95.625 94.065 ;
        RECT 93.375 93.410 94.595 93.425 ;
        RECT 63.830 92.635 66.340 92.935 ;
        RECT 54.715 83.090 55.845 83.525 ;
        RECT 53.465 82.790 55.845 83.090 ;
        RECT 52.285 76.945 53.015 77.180 ;
        RECT 53.465 76.945 53.765 82.790 ;
        RECT 54.715 82.355 55.845 82.790 ;
        RECT 63.830 83.185 64.130 92.635 ;
        RECT 65.210 92.325 66.340 92.635 ;
        RECT 91.330 92.710 94.595 93.410 ;
        RECT 104.530 93.135 105.660 94.305 ;
        RECT 111.790 94.065 113.955 94.765 ;
        RECT 111.790 93.495 112.490 94.065 ;
        RECT 112.825 93.820 113.955 94.065 ;
        RECT 109.660 93.425 112.710 93.495 ;
        RECT 91.330 91.920 92.030 92.710 ;
        RECT 93.465 92.255 94.595 92.710 ;
        RECT 109.660 92.795 112.925 93.425 ;
        RECT 109.660 91.920 110.360 92.795 ;
        RECT 111.795 92.255 112.925 92.795 ;
        RECT 91.115 91.540 92.245 91.920 ;
        RECT 109.445 91.625 110.575 91.920 ;
        RECT 88.160 90.840 92.245 91.540 ;
        RECT 88.160 89.760 88.860 90.840 ;
        RECT 91.115 90.750 92.245 90.840 ;
        RECT 106.490 90.925 110.575 91.625 ;
        RECT 106.490 89.780 107.190 90.925 ;
        RECT 109.445 90.750 110.575 90.925 ;
        RECT 87.900 88.590 89.030 89.760 ;
        RECT 106.230 88.610 107.360 89.780 ;
        RECT 88.175 87.005 88.875 88.590 ;
        RECT 90.435 87.005 91.565 87.380 ;
        RECT 88.175 86.305 91.565 87.005 ;
        RECT 106.505 87.145 107.205 88.610 ;
        RECT 108.765 87.145 109.895 87.380 ;
        RECT 106.505 86.445 109.895 87.145 ;
        RECT 90.435 86.210 91.565 86.305 ;
        RECT 108.765 86.210 109.895 86.445 ;
        RECT 90.790 85.230 91.490 86.210 ;
        RECT 92.510 85.230 93.640 85.955 ;
        RECT 90.790 84.785 93.640 85.230 ;
        RECT 109.120 85.370 109.820 86.210 ;
        RECT 110.840 85.370 111.970 85.955 ;
        RECT 109.120 84.785 111.970 85.370 ;
        RECT 90.790 84.530 93.425 84.785 ;
        RECT 109.120 84.670 111.755 84.785 ;
        RECT 92.725 84.010 93.425 84.530 ;
        RECT 111.055 84.010 111.755 84.670 ;
        RECT 65.210 83.185 66.340 83.640 ;
        RECT 74.255 83.390 75.385 83.790 ;
        RECT 63.830 82.885 66.340 83.185 ;
        RECT 52.285 76.645 53.765 76.945 ;
        RECT 52.285 76.410 53.015 76.645 ;
        RECT 45.730 73.910 46.860 74.345 ;
        RECT 53.465 74.210 53.765 76.645 ;
        RECT 54.715 74.220 55.845 74.320 ;
        RECT 63.830 74.220 64.130 82.885 ;
        RECT 65.210 82.470 66.340 82.885 ;
        RECT 72.705 83.090 75.385 83.390 ;
        RECT 65.210 74.220 66.340 74.465 ;
        RECT 54.715 74.210 66.340 74.220 ;
        RECT 53.465 73.920 66.340 74.210 ;
        RECT 53.465 73.910 55.845 73.920 ;
        RECT 45.730 73.790 53.765 73.910 ;
        RECT 44.765 73.610 53.765 73.790 ;
        RECT 44.765 73.490 46.860 73.610 ;
        RECT 45.730 73.175 46.860 73.490 ;
        RECT 54.715 73.150 55.845 73.910 ;
        RECT 65.210 73.295 66.340 73.920 ;
        RECT 72.705 73.700 73.005 83.090 ;
        RECT 74.255 82.620 75.385 83.090 ;
        RECT 92.510 82.840 93.640 84.010 ;
        RECT 110.840 82.840 111.970 84.010 ;
        RECT 92.590 82.095 93.290 82.840 ;
        RECT 94.780 82.095 95.910 82.470 ;
        RECT 92.590 81.395 95.910 82.095 ;
        RECT 94.780 81.300 95.910 81.395 ;
        RECT 97.935 82.115 99.065 82.470 ;
        RECT 110.920 82.115 111.620 82.840 ;
        RECT 113.110 82.115 114.240 82.470 ;
        RECT 97.935 81.415 114.240 82.115 ;
        RECT 97.935 81.300 99.065 81.415 ;
        RECT 94.995 80.975 95.695 81.300 ;
        RECT 98.160 80.975 98.860 81.300 ;
        RECT 94.995 80.275 98.860 80.975 ;
        RECT 96.160 78.230 97.290 78.425 ;
        RECT 94.420 77.530 97.290 78.230 ;
        RECT 94.420 76.700 95.120 77.530 ;
        RECT 96.160 77.255 97.290 77.530 ;
        RECT 94.205 76.475 95.335 76.700 ;
        RECT 93.190 75.775 95.335 76.475 ;
        RECT 93.190 75.265 93.890 75.775 ;
        RECT 94.205 75.530 95.335 75.775 ;
        RECT 90.845 75.135 93.895 75.265 ;
        RECT 90.845 74.565 94.305 75.135 ;
        RECT 73.850 73.700 74.980 74.165 ;
        RECT 72.705 73.400 74.980 73.700 ;
        RECT 90.845 73.630 91.545 74.565 ;
        RECT 93.175 73.965 94.305 74.565 ;
        RECT 72.705 72.850 73.005 73.400 ;
        RECT 73.850 72.995 74.980 73.400 ;
        RECT 90.825 73.395 91.955 73.630 ;
        RECT 50.435 72.550 73.005 72.850 ;
        RECT 87.675 72.695 91.955 73.395 ;
        RECT 50.435 66.710 50.735 72.550 ;
        RECT 58.390 70.285 58.690 72.550 ;
        RECT 87.675 71.490 88.375 72.695 ;
        RECT 90.825 72.460 91.955 72.695 ;
        RECT 87.610 70.320 88.740 71.490 ;
        RECT 58.205 69.515 58.935 70.285 ;
        RECT 87.675 68.625 88.375 70.320 ;
        RECT 90.145 68.625 91.275 69.090 ;
        RECT 87.675 67.925 91.275 68.625 ;
        RECT 90.145 67.920 91.275 67.925 ;
        RECT 51.325 66.710 52.455 67.145 ;
        RECT 50.435 66.410 52.455 66.710 ;
        RECT 47.765 59.970 48.495 60.250 ;
        RECT 50.435 59.970 50.735 66.410 ;
        RECT 51.325 65.975 52.455 66.410 ;
        RECT 90.500 66.850 91.200 67.920 ;
        RECT 92.220 66.850 93.350 67.665 ;
        RECT 90.500 66.495 93.350 66.850 ;
        RECT 90.500 66.150 93.135 66.495 ;
        RECT 92.435 65.720 93.135 66.150 ;
        RECT 92.220 64.550 93.350 65.720 ;
        RECT 92.300 63.715 93.000 64.550 ;
        RECT 94.490 63.715 95.620 64.180 ;
        RECT 92.300 63.015 95.620 63.715 ;
        RECT 94.490 63.010 95.620 63.015 ;
        RECT 97.645 63.480 98.775 64.180 ;
        RECT 103.265 63.480 103.965 81.415 ;
        RECT 113.110 81.300 114.240 81.415 ;
        RECT 116.265 81.300 117.395 82.470 ;
        RECT 113.455 80.995 114.155 81.300 ;
        RECT 116.480 80.995 117.180 81.300 ;
        RECT 113.455 80.295 117.180 80.995 ;
        RECT 114.760 77.985 115.890 78.180 ;
        RECT 113.070 77.285 115.890 77.985 ;
        RECT 113.070 76.455 113.770 77.285 ;
        RECT 114.760 77.010 115.890 77.285 ;
        RECT 112.855 76.230 113.985 76.455 ;
        RECT 111.815 75.530 113.985 76.230 ;
        RECT 111.815 75.020 112.515 75.530 ;
        RECT 112.855 75.285 113.985 75.530 ;
        RECT 109.475 74.890 112.525 75.020 ;
        RECT 109.475 74.320 112.955 74.890 ;
        RECT 109.475 73.385 110.175 74.320 ;
        RECT 111.815 74.305 112.955 74.320 ;
        RECT 111.825 73.720 112.955 74.305 ;
        RECT 109.475 73.150 110.605 73.385 ;
        RECT 106.305 72.450 110.605 73.150 ;
        RECT 106.305 71.260 107.005 72.450 ;
        RECT 109.475 72.215 110.605 72.450 ;
        RECT 106.260 70.090 107.390 71.260 ;
        RECT 106.305 68.610 107.005 70.090 ;
        RECT 108.795 68.610 109.925 68.845 ;
        RECT 106.305 67.910 109.925 68.610 ;
        RECT 108.795 67.675 109.925 67.910 ;
        RECT 109.150 66.835 109.850 67.675 ;
        RECT 110.870 66.835 112.000 67.420 ;
        RECT 109.150 66.250 112.000 66.835 ;
        RECT 109.150 66.135 111.785 66.250 ;
        RECT 111.085 65.475 111.785 66.135 ;
        RECT 110.870 64.305 112.000 65.475 ;
        RECT 110.950 63.480 111.650 64.305 ;
        RECT 113.140 63.480 114.270 63.935 ;
        RECT 97.645 63.010 114.270 63.480 ;
        RECT 94.705 62.595 95.405 63.010 ;
        RECT 97.860 62.780 114.270 63.010 ;
        RECT 97.860 62.595 98.570 62.780 ;
        RECT 94.705 61.895 98.570 62.595 ;
        RECT 102.375 62.115 103.075 62.780 ;
        RECT 113.140 62.765 114.270 62.780 ;
        RECT 116.295 62.765 117.425 63.935 ;
        RECT 113.355 62.360 114.055 62.765 ;
        RECT 116.520 62.360 117.220 62.765 ;
        RECT 102.375 61.375 103.150 62.115 ;
        RECT 113.355 61.660 117.220 62.360 ;
        RECT 102.430 61.335 103.150 61.375 ;
        RECT 51.325 59.970 52.455 60.455 ;
        RECT 47.765 59.670 52.455 59.970 ;
        RECT 47.765 59.480 48.495 59.670 ;
        RECT 51.325 59.285 52.455 59.670 ;
        RECT 105.140 60.085 109.810 60.115 ;
        RECT 105.140 59.415 112.410 60.085 ;
        RECT 105.140 56.670 105.840 59.415 ;
        RECT 108.730 59.385 112.410 59.415 ;
        RECT 108.730 58.300 109.430 59.385 ;
        RECT 111.710 58.300 112.410 59.385 ;
        RECT 108.495 57.130 109.625 58.300 ;
        RECT 111.495 57.130 112.625 58.300 ;
        RECT 106.245 56.670 107.375 56.890 ;
        RECT 72.780 55.325 73.900 56.505 ;
        RECT 103.945 55.970 107.375 56.670 ;
        RECT 103.945 54.780 104.645 55.970 ;
        RECT 106.245 55.720 107.375 55.970 ;
        RECT 105.910 54.780 107.040 55.215 ;
        RECT 103.945 54.480 107.040 54.780 ;
        RECT 51.325 53.355 52.455 53.790 ;
        RECT 50.425 53.055 52.455 53.355 ;
        RECT 50.425 46.875 50.725 53.055 ;
        RECT 51.325 52.620 52.455 53.055 ;
        RECT 61.340 50.730 62.470 51.900 ;
        RECT 72.780 51.575 73.900 52.755 ;
        RECT 103.945 51.740 104.645 54.480 ;
        RECT 105.910 54.045 107.040 54.480 ;
        RECT 103.945 51.160 104.710 51.740 ;
        RECT 105.910 51.160 107.040 51.595 ;
        RECT 103.945 51.040 107.040 51.160 ;
        RECT 59.825 49.405 60.955 50.575 ;
        RECT 61.755 50.015 62.055 50.730 ;
        RECT 60.365 47.860 60.665 49.405 ;
        RECT 61.340 48.845 62.470 50.015 ;
        RECT 72.875 49.845 74.005 51.015 ;
        RECT 104.005 50.860 107.040 51.040 ;
        RECT 61.755 48.190 62.055 48.845 ;
        RECT 73.340 48.445 73.640 49.845 ;
        RECT 61.340 47.860 62.470 48.190 ;
        RECT 60.365 47.560 62.470 47.860 ;
        RECT 51.325 46.965 52.455 47.165 ;
        RECT 60.365 46.965 60.665 47.560 ;
        RECT 61.340 47.020 62.470 47.560 ;
        RECT 72.815 47.275 73.945 48.445 ;
        RECT 51.325 46.875 60.665 46.965 ;
        RECT 50.425 46.665 60.665 46.875 ;
        RECT 50.425 46.575 52.455 46.665 ;
        RECT 51.325 45.995 52.455 46.575 ;
        RECT 61.755 46.315 62.055 47.020 ;
        RECT 61.340 45.145 62.470 46.315 ;
        RECT 73.340 45.940 73.640 47.275 ;
        RECT 104.005 46.005 104.705 50.860 ;
        RECT 105.910 50.425 107.040 50.860 ;
        RECT 105.910 47.610 107.040 47.845 ;
        RECT 105.565 46.675 107.040 47.610 ;
        RECT 105.565 46.005 106.265 46.675 ;
        RECT 106.585 46.005 107.715 46.240 ;
        RECT 61.755 44.495 62.055 45.145 ;
        RECT 72.925 44.770 74.055 45.940 ;
        RECT 104.005 45.305 107.715 46.005 ;
        RECT 61.340 43.325 62.470 44.495 ;
        RECT 73.340 43.330 73.640 44.770 ;
        RECT 61.755 42.755 62.055 43.325 ;
        RECT 61.340 41.585 62.470 42.755 ;
        RECT 72.925 42.160 74.055 43.330 ;
        RECT 36.860 40.500 38.500 40.530 ;
        RECT 39.250 40.500 40.380 40.935 ;
        RECT 48.060 40.510 49.190 40.945 ;
        RECT 61.755 40.920 62.055 41.585 ;
        RECT 36.860 40.200 40.380 40.500 ;
        RECT 36.860 34.030 37.160 40.200 ;
        RECT 39.250 39.765 40.380 40.200 ;
        RECT 45.885 40.210 49.190 40.510 ;
        RECT 38.900 34.030 40.030 34.230 ;
        RECT 36.860 33.730 40.030 34.030 ;
        RECT 36.860 27.810 37.160 33.730 ;
        RECT 38.900 33.060 40.030 33.730 ;
        RECT 45.885 33.815 46.185 40.210 ;
        RECT 48.060 39.775 49.190 40.210 ;
        RECT 61.340 39.750 62.470 40.920 ;
        RECT 73.340 40.845 73.640 42.160 ;
        RECT 97.120 41.740 98.250 42.230 ;
        RECT 105.565 41.740 106.265 45.305 ;
        RECT 106.585 45.070 107.715 45.305 ;
        RECT 108.995 43.580 110.125 44.750 ;
        RECT 111.725 43.620 112.855 44.790 ;
        RECT 109.240 41.740 109.940 43.580 ;
        RECT 111.940 41.740 112.640 43.620 ;
        RECT 97.120 41.060 112.640 41.740 ;
        RECT 97.335 41.040 112.640 41.060 ;
        RECT 72.925 39.675 74.055 40.845 ;
        RECT 73.340 38.960 73.640 39.675 ;
        RECT 73.010 38.190 73.740 38.960 ;
        RECT 58.900 36.275 60.030 36.710 ;
        RECT 72.740 36.275 73.870 37.070 ;
        RECT 56.085 35.975 73.870 36.275 ;
        RECT 48.045 33.870 49.175 34.240 ;
        RECT 56.085 33.870 56.385 35.975 ;
        RECT 58.900 35.540 60.030 35.975 ;
        RECT 72.740 35.900 73.870 35.975 ;
        RECT 45.885 33.805 47.070 33.815 ;
        RECT 48.045 33.805 56.385 33.870 ;
        RECT 45.885 33.570 56.385 33.805 ;
        RECT 45.885 33.505 49.175 33.570 ;
        RECT 38.900 27.810 40.030 28.115 ;
        RECT 36.860 27.510 40.030 27.810 ;
        RECT 36.860 21.285 37.160 27.510 ;
        RECT 38.900 26.945 40.030 27.510 ;
        RECT 45.885 27.780 46.185 33.505 ;
        RECT 48.045 33.070 49.175 33.505 ;
        RECT 57.715 33.230 58.435 33.355 ;
        RECT 58.900 33.230 60.030 33.665 ;
        RECT 57.715 32.930 60.030 33.230 ;
        RECT 57.715 32.575 58.435 32.930 ;
        RECT 58.900 32.495 60.030 32.930 ;
        RECT 48.080 27.780 49.210 28.145 ;
        RECT 45.885 27.480 49.210 27.780 ;
        RECT 37.910 21.285 39.040 21.720 ;
        RECT 36.860 21.200 39.040 21.285 ;
        RECT 45.885 21.200 46.185 27.480 ;
        RECT 46.815 27.460 47.115 27.480 ;
        RECT 48.080 26.975 49.210 27.480 ;
        RECT 48.035 21.200 49.165 21.740 ;
        RECT 36.860 20.985 49.165 21.200 ;
        RECT 37.910 20.900 49.165 20.985 ;
        RECT 37.910 20.550 39.040 20.900 ;
        RECT 48.035 20.570 49.165 20.900 ;
        RECT 97.120 19.435 98.250 19.870 ;
        RECT 102.050 19.435 124.505 35.935 ;
        RECT 97.120 19.135 124.505 19.435 ;
        RECT 97.120 18.700 98.250 19.135 ;
        RECT 102.050 13.485 124.505 19.135 ;
        RECT 134.200 4.555 135.370 4.560 ;
        RECT 154.755 4.555 155.925 4.560 ;
        RECT 112.225 4.215 113.395 4.220 ;
        RECT 112.220 3.095 113.400 4.215 ;
        RECT 134.195 3.435 135.375 4.555 ;
        RECT 154.750 3.435 155.930 4.555 ;
        RECT 134.200 3.430 135.370 3.435 ;
        RECT 154.755 3.430 155.925 3.435 ;
        RECT 112.225 3.090 113.395 3.095 ;
      LAYER met4 ;
        RECT 3.490 225.040 3.990 225.055 ;
        RECT 4.290 225.040 7.670 225.055 ;
        RECT 5.490 224.760 7.670 225.040 ;
        RECT 7.970 224.760 11.350 225.055 ;
        RECT 11.650 224.760 15.030 225.055 ;
        RECT 15.330 224.760 18.710 225.055 ;
        RECT 19.010 224.760 22.390 225.055 ;
        RECT 22.690 224.760 26.070 225.055 ;
        RECT 26.370 224.760 29.750 225.055 ;
        RECT 30.050 224.760 33.430 225.055 ;
        RECT 33.730 224.760 37.110 225.055 ;
        RECT 37.410 224.760 40.790 225.055 ;
        RECT 41.090 224.760 44.470 225.055 ;
        RECT 44.770 224.760 48.150 225.055 ;
        RECT 48.450 224.760 51.830 225.055 ;
        RECT 52.130 224.760 55.510 225.055 ;
        RECT 55.810 224.760 59.190 225.055 ;
        RECT 59.490 224.760 62.870 225.055 ;
        RECT 63.170 224.760 66.550 225.055 ;
        RECT 66.850 224.760 70.230 225.055 ;
        RECT 70.530 224.760 73.910 225.055 ;
        RECT 74.210 224.760 77.590 225.055 ;
        RECT 77.890 224.760 81.270 225.055 ;
        RECT 81.570 224.760 84.950 225.055 ;
        RECT 85.250 224.760 88.630 225.055 ;
        RECT 5.490 224.755 88.770 224.760 ;
        RECT 158.355 224.145 160.355 224.150 ;
        RECT 56.955 219.580 58.085 219.645 ;
        RECT 15.025 218.580 58.085 219.580 ;
        RECT 7.815 214.665 8.945 214.730 ;
        RECT 5.490 213.665 8.945 214.665 ;
        RECT 7.815 213.600 8.945 213.665 ;
        RECT 7.815 110.755 8.945 110.820 ;
        RECT 5.490 109.755 8.945 110.755 ;
        RECT 7.815 109.690 8.945 109.755 ;
        RECT 15.025 2.675 16.025 218.580 ;
        RECT 56.955 218.515 58.085 218.580 ;
        RECT 132.115 215.925 133.245 215.990 ;
        RECT 158.355 215.925 158.360 224.145 ;
        RECT 132.115 214.925 158.360 215.925 ;
        RECT 132.115 214.860 133.245 214.925 ;
        RECT 111.315 123.660 112.445 123.725 ;
        RECT 20.500 122.660 112.445 123.660 ;
        RECT 20.500 4.570 21.500 122.660 ;
        RECT 111.315 122.595 112.445 122.660 ;
        RECT 137.770 110.335 138.900 110.400 ;
        RECT 158.355 110.335 158.360 214.925 ;
        RECT 137.770 109.335 158.360 110.335 ;
        RECT 137.770 109.270 138.900 109.335 ;
        RECT 102.425 61.360 103.155 62.090 ;
        RECT 72.775 55.350 73.905 56.480 ;
        RECT 73.190 53.445 73.490 55.350 ;
        RECT 59.390 53.145 73.490 53.445 ;
        RECT 59.390 44.920 59.690 53.145 ;
        RECT 73.190 52.730 73.490 53.145 ;
        RECT 72.775 51.600 73.905 52.730 ;
        RECT 57.770 44.900 59.690 44.920 ;
        RECT 56.755 44.620 59.690 44.900 ;
        RECT 56.755 44.600 58.070 44.620 ;
        RECT 56.755 33.115 57.055 44.600 ;
        RECT 102.440 35.795 103.140 61.360 ;
        RECT 57.710 33.115 58.440 33.330 ;
        RECT 56.755 32.815 58.440 33.115 ;
        RECT 57.710 32.600 58.440 32.815 ;
        RECT 102.190 13.625 124.365 35.795 ;
        RECT 90.070 4.570 91.160 4.600 ;
        RECT 20.500 3.570 91.160 4.570 ;
        RECT 15.025 1.675 69.045 2.675 ;
        RECT 68.045 1.000 69.045 1.675 ;
        RECT 68.045 0.495 68.090 1.000 ;
        RECT 68.990 0.495 69.045 1.000 ;
        RECT 90.070 1.000 91.160 3.570 ;
        RECT 112.245 3.380 113.375 4.220 ;
        RECT 134.220 3.430 135.350 4.560 ;
        RECT 154.775 4.495 155.905 4.560 ;
        RECT 154.775 3.495 157.405 4.495 ;
        RECT 154.775 3.430 155.905 3.495 ;
        RECT 90.070 0.470 90.170 1.000 ;
        RECT 91.070 0.470 91.160 1.000 ;
        RECT 112.090 1.000 113.390 3.380 ;
        RECT 112.090 0.530 112.250 1.000 ;
        RECT 113.150 0.530 113.390 1.000 ;
        RECT 134.285 1.000 135.285 3.430 ;
        RECT 134.285 0.460 134.330 1.000 ;
        RECT 135.230 0.460 135.285 1.000 ;
        RECT 156.340 1.000 157.405 3.495 ;
        RECT 156.340 0.460 156.410 1.000 ;
        RECT 157.310 0.470 157.405 1.000 ;
        RECT 157.310 0.460 157.400 0.470 ;
        RECT 158.355 0.265 158.360 109.335 ;
  END
END tt_um_Burrows_Katie
END LIBRARY

