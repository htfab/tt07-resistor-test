VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Burrows_Katie
  CLASS BLOCK ;
  FOREIGN tt_um_Burrows_Katie ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.860 225.760 155.160 225.770 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.540 225.760 158.840 225.770 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.980 225.760 4.280 225.770 ;
        RECT 7.660 225.760 7.960 225.770 ;
        RECT 11.340 225.760 11.640 225.770 ;
        RECT 15.020 225.760 15.320 225.770 ;
        RECT 18.700 225.760 19.000 225.770 ;
        RECT 22.380 225.760 22.680 225.770 ;
        RECT 26.060 225.760 26.360 225.770 ;
        RECT 29.740 225.760 30.040 225.770 ;
        RECT 33.420 225.760 33.720 225.770 ;
        RECT 37.100 225.760 37.400 225.770 ;
        RECT 40.780 225.760 41.080 225.770 ;
        RECT 44.460 225.760 44.760 225.770 ;
        RECT 48.140 225.760 48.440 225.770 ;
        RECT 51.820 225.760 52.120 225.770 ;
        RECT 55.500 225.760 55.800 225.770 ;
        RECT 59.180 225.760 59.480 225.770 ;
        RECT 62.860 225.760 63.160 225.770 ;
        RECT 66.540 225.760 66.840 225.770 ;
        RECT 70.220 225.760 70.520 225.770 ;
        RECT 73.900 225.760 74.200 225.770 ;
        RECT 77.580 225.760 77.880 225.770 ;
        RECT 81.260 225.760 81.560 225.770 ;
        RECT 84.940 225.760 85.240 225.770 ;
        RECT 88.620 225.760 88.920 225.770 ;
        RECT 4.585 54.895 4.595 54.905 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.180 225.760 151.480 225.770 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.280 43.405 159.290 43.415 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 17.639999 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.410000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.410000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.095000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.500 225.760 147.800 225.770 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.820 225.760 144.120 225.770 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.140 225.760 140.440 225.770 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.460 225.760 136.760 225.770 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.780 225.760 133.080 225.770 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.100 225.760 129.400 225.770 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.420 225.760 125.720 225.770 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.740 225.760 122.040 225.770 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.060 225.760 118.360 225.770 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.380 225.760 114.680 225.770 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.700 225.760 111.000 225.770 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.020 225.760 107.320 225.770 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.340 225.760 103.640 225.770 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.660 225.760 99.960 225.770 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.980 225.760 96.280 225.770 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.300 225.760 92.600 225.770 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 78.979797 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER pwell ;
        RECT 52.635 212.190 53.305 212.270 ;
        RECT 52.635 209.400 58.575 212.190 ;
      LAYER nwell ;
        RECT 98.110 210.380 104.530 215.660 ;
        RECT 106.190 210.380 112.610 215.660 ;
      LAYER pwell ;
        RECT 52.635 209.320 53.305 209.400 ;
        RECT 52.635 207.490 53.305 207.570 ;
        RECT 52.635 204.700 58.575 207.490 ;
      LAYER nwell ;
        RECT 63.295 206.310 65.715 209.590 ;
        RECT 92.275 206.345 94.695 209.625 ;
      LAYER pwell ;
        RECT 52.635 204.620 53.305 204.700 ;
      LAYER nwell ;
        RECT 98.110 203.390 104.530 208.670 ;
        RECT 106.190 203.390 112.610 208.670 ;
      LAYER pwell ;
        RECT 52.635 200.955 53.305 201.035 ;
        RECT 52.635 198.165 58.575 200.955 ;
        RECT 52.635 198.085 53.305 198.165 ;
      LAYER nwell ;
        RECT 76.820 197.000 83.240 202.280 ;
        RECT 98.110 196.400 104.530 201.680 ;
        RECT 106.190 196.400 112.610 201.680 ;
      LAYER pwell ;
        RECT 52.635 196.145 53.305 196.225 ;
        RECT 52.635 193.355 58.575 196.145 ;
        RECT 52.635 193.275 53.305 193.355 ;
      LAYER nwell ;
        RECT 76.820 190.085 83.240 195.365 ;
        RECT 98.110 189.375 104.530 194.655 ;
        RECT 106.190 189.375 112.610 194.655 ;
      LAYER pwell ;
        RECT 45.540 187.750 46.210 187.830 ;
        RECT 45.540 184.960 53.480 187.750 ;
        RECT 45.540 184.880 46.210 184.960 ;
        RECT 45.540 183.275 46.210 183.355 ;
        RECT 45.540 180.485 53.480 183.275 ;
        RECT 45.540 180.405 46.210 180.485 ;
        RECT 45.540 178.660 46.210 178.740 ;
        RECT 45.540 175.870 53.480 178.660 ;
        RECT 45.540 175.790 46.210 175.870 ;
        RECT 45.520 173.085 46.190 173.165 ;
        RECT 45.520 170.295 53.460 173.085 ;
      LAYER nwell ;
        RECT 88.670 172.375 91.090 175.655 ;
        RECT 106.415 170.760 112.835 176.040 ;
      LAYER pwell ;
        RECT 45.520 170.215 46.190 170.295 ;
        RECT 45.520 168.570 46.190 168.650 ;
        RECT 45.520 165.780 53.460 168.570 ;
        RECT 45.520 165.700 46.190 165.780 ;
        RECT 45.520 163.980 46.190 164.060 ;
        RECT 45.520 161.190 53.460 163.980 ;
      LAYER nwell ;
        RECT 88.665 162.375 91.085 165.655 ;
        RECT 106.415 163.650 112.835 168.930 ;
      LAYER pwell ;
        RECT 45.520 161.110 46.190 161.190 ;
        RECT 43.420 107.235 44.090 107.315 ;
        RECT 43.420 102.445 49.360 107.235 ;
        RECT 43.420 102.365 44.090 102.445 ;
      LAYER nwell ;
        RECT 52.685 102.255 59.105 107.535 ;
        RECT 62.835 102.255 69.255 107.535 ;
        RECT 72.115 102.210 78.535 107.490 ;
      LAYER pwell ;
        RECT 43.420 97.420 44.090 97.500 ;
        RECT 43.420 92.630 49.360 97.420 ;
        RECT 43.420 92.550 44.090 92.630 ;
      LAYER nwell ;
        RECT 52.685 92.360 59.105 97.640 ;
        RECT 62.835 92.380 69.255 97.660 ;
        RECT 72.115 92.320 78.535 97.600 ;
      LAYER pwell ;
        RECT 43.420 87.260 44.090 87.340 ;
        RECT 43.420 82.470 49.360 87.260 ;
        RECT 43.420 82.390 44.090 82.470 ;
      LAYER nwell ;
        RECT 52.685 82.315 59.105 87.595 ;
        RECT 62.835 82.440 69.255 87.720 ;
        RECT 72.070 82.485 78.490 87.765 ;
        RECT 95.515 81.225 101.935 94.195 ;
        RECT 113.860 81.225 120.280 94.195 ;
      LAYER pwell ;
        RECT 43.420 78.195 44.090 78.275 ;
        RECT 43.420 73.405 49.360 78.195 ;
        RECT 43.420 73.325 44.090 73.405 ;
      LAYER nwell ;
        RECT 52.685 73.115 59.105 78.395 ;
        RECT 62.835 73.020 69.255 78.300 ;
        RECT 72.115 72.925 78.535 78.205 ;
      LAYER pwell ;
        RECT 49.105 69.980 49.775 70.060 ;
        RECT 49.105 66.190 56.045 69.980 ;
        RECT 49.105 66.110 49.775 66.190 ;
        RECT 49.105 63.290 49.775 63.370 ;
        RECT 49.105 59.500 56.045 63.290 ;
        RECT 49.105 59.420 49.775 59.500 ;
        RECT 49.105 56.600 49.775 56.680 ;
        RECT 49.105 52.810 56.045 56.600 ;
      LAYER nwell ;
        RECT 62.030 54.460 70.450 68.200 ;
        RECT 74.385 54.880 82.805 68.680 ;
        RECT 95.210 62.935 101.630 75.905 ;
        RECT 113.865 62.690 120.285 75.660 ;
      LAYER pwell ;
        RECT 49.105 52.730 49.775 52.810 ;
        RECT 49.105 49.960 49.775 50.040 ;
        RECT 49.105 46.170 56.045 49.960 ;
        RECT 49.105 46.090 49.775 46.170 ;
        RECT 35.635 43.760 36.305 43.840 ;
        RECT 45.760 43.760 46.430 43.840 ;
        RECT 35.635 39.970 42.675 43.760 ;
        RECT 45.760 39.970 52.800 43.760 ;
        RECT 35.635 39.890 36.305 39.970 ;
        RECT 45.760 39.890 46.430 39.970 ;
      LAYER nwell ;
        RECT 62.285 37.755 70.705 51.495 ;
        RECT 74.405 37.235 82.825 51.035 ;
        RECT 111.050 43.660 119.470 56.000 ;
      LAYER pwell ;
        RECT 35.635 37.065 36.305 37.145 ;
        RECT 45.760 37.065 46.430 37.145 ;
        RECT 35.635 33.275 42.675 37.065 ;
        RECT 45.760 33.275 52.800 37.065 ;
        RECT 70.115 34.305 70.785 34.385 ;
        RECT 56.665 34.130 57.335 34.210 ;
        RECT 35.635 33.195 36.305 33.275 ;
        RECT 45.760 33.195 46.430 33.275 ;
        RECT 56.665 32.710 64.605 34.130 ;
        RECT 70.115 32.885 78.055 34.305 ;
        RECT 70.115 32.805 70.785 32.885 ;
        RECT 56.665 32.630 57.335 32.710 ;
        RECT 35.635 30.950 36.305 31.030 ;
        RECT 45.760 30.950 46.430 31.030 ;
        RECT 35.635 27.160 42.675 30.950 ;
        RECT 45.760 27.160 52.800 30.950 ;
        RECT 35.635 27.080 36.305 27.160 ;
        RECT 45.760 27.080 46.430 27.160 ;
        RECT 35.635 24.545 36.305 24.625 ;
        RECT 45.760 24.545 46.430 24.625 ;
        RECT 35.635 20.755 42.675 24.545 ;
        RECT 45.760 20.755 52.800 24.545 ;
        RECT 35.635 20.675 36.305 20.755 ;
        RECT 45.760 20.675 46.430 20.755 ;
      LAYER li1 ;
        RECT 98.985 215.640 99.515 216.170 ;
        RECT 107.265 215.640 107.795 216.170 ;
        RECT 99.100 215.245 99.400 215.640 ;
        RECT 98.795 215.075 103.545 215.245 ;
        RECT 103.980 214.580 104.310 215.325 ;
        RECT 107.380 215.245 107.680 215.640 ;
        RECT 106.875 215.075 111.625 215.245 ;
        RECT 104.595 214.580 105.125 214.715 ;
        RECT 103.980 214.250 105.125 214.580 ;
        RECT 52.805 211.275 53.135 212.100 ;
        RECT 53.840 212.020 54.540 213.210 ;
        RECT 97.590 212.980 98.190 213.580 ;
        RECT 53.570 211.850 58.320 212.020 ;
        RECT 51.895 210.575 53.135 211.275 ;
        RECT 52.805 209.490 53.135 210.575 ;
        RECT 59.000 210.430 59.530 210.960 ;
        RECT 98.795 210.795 103.545 210.965 ;
        RECT 103.230 210.380 103.400 210.795 ;
        RECT 103.980 210.715 104.310 214.250 ;
        RECT 104.595 214.185 105.125 214.250 ;
        RECT 112.060 214.425 112.390 215.325 ;
        RECT 112.695 214.425 113.225 214.565 ;
        RECT 112.060 214.095 113.225 214.425 ;
        RECT 105.785 213.120 106.385 213.720 ;
        RECT 106.875 210.795 111.625 210.965 ;
        RECT 107.080 210.650 107.385 210.795 ;
        RECT 112.060 210.715 112.390 214.095 ;
        RECT 112.695 214.035 113.225 214.095 ;
        RECT 107.085 210.380 107.385 210.650 ;
        RECT 53.570 209.570 58.320 209.740 ;
        RECT 64.100 209.640 64.630 210.170 ;
        RECT 93.185 209.640 93.715 210.170 ;
        RECT 103.050 209.850 103.580 210.380 ;
        RECT 106.970 209.850 107.500 210.380 ;
        RECT 53.640 209.240 53.940 209.570 ;
        RECT 53.525 208.710 54.055 209.240 ;
        RECT 64.215 209.175 64.385 209.640 ;
        RECT 65.185 209.255 65.515 209.275 ;
        RECT 64.020 209.005 64.690 209.175 ;
        RECT 52.805 206.375 53.135 207.400 ;
        RECT 53.830 207.320 54.530 208.145 ;
        RECT 62.560 207.930 63.450 208.820 ;
        RECT 53.570 207.150 58.320 207.320 ;
        RECT 64.020 206.830 64.690 206.895 ;
        RECT 51.895 205.675 53.135 206.375 ;
        RECT 64.005 206.725 64.690 206.830 ;
        RECT 64.005 206.365 64.405 206.725 ;
        RECT 65.165 206.645 65.515 209.255 ;
        RECT 93.310 209.210 93.610 209.640 ;
        RECT 93.000 209.040 93.670 209.210 ;
        RECT 93.310 209.005 93.610 209.040 ;
        RECT 91.470 207.930 92.360 208.820 ;
        RECT 93.000 206.760 93.670 206.930 ;
        RECT 94.145 206.820 94.475 209.290 ;
        RECT 98.985 208.445 99.515 208.975 ;
        RECT 107.265 208.445 107.795 208.975 ;
        RECT 99.100 208.255 99.400 208.445 ;
        RECT 98.795 208.085 103.545 208.255 ;
        RECT 59.000 205.775 59.530 206.305 ;
        RECT 63.920 205.835 64.450 206.365 ;
        RECT 52.805 204.790 53.135 205.675 ;
        RECT 65.185 205.290 65.515 206.645 ;
        RECT 93.310 206.385 93.610 206.760 ;
        RECT 94.120 206.680 94.475 206.820 ;
        RECT 103.980 207.660 104.310 208.335 ;
        RECT 107.380 208.255 107.680 208.445 ;
        RECT 106.875 208.085 111.625 208.255 ;
        RECT 104.615 207.660 105.145 207.800 ;
        RECT 103.980 207.330 105.145 207.660 ;
        RECT 93.185 205.855 93.715 206.385 ;
        RECT 94.120 205.385 94.450 206.680 ;
        RECT 97.590 205.805 98.190 206.405 ;
        RECT 53.570 204.870 58.320 205.040 ;
        RECT 53.600 204.430 53.900 204.870 ;
        RECT 65.185 204.860 65.725 205.290 ;
        RECT 65.195 204.760 65.725 204.860 ;
        RECT 93.995 204.855 94.525 205.385 ;
        RECT 53.485 203.900 54.015 204.430 ;
        RECT 98.795 203.805 103.545 203.975 ;
        RECT 103.315 203.315 103.485 203.805 ;
        RECT 103.980 203.725 104.310 207.330 ;
        RECT 104.615 207.270 105.145 207.330 ;
        RECT 112.060 207.660 112.390 208.335 ;
        RECT 112.695 207.660 113.225 207.800 ;
        RECT 112.060 207.330 113.225 207.660 ;
        RECT 105.785 206.040 106.385 206.640 ;
        RECT 106.875 203.805 111.625 203.975 ;
        RECT 107.170 203.315 107.470 203.805 ;
        RECT 112.060 203.725 112.390 207.330 ;
        RECT 112.695 207.270 113.225 207.330 ;
        RECT 81.465 201.865 82.165 203.085 ;
        RECT 103.135 202.785 103.665 203.315 ;
        RECT 107.055 202.785 107.585 203.315 ;
        RECT 52.805 199.840 53.135 200.865 ;
        RECT 53.755 200.785 54.455 201.715 ;
        RECT 77.505 201.695 82.255 201.865 ;
        RECT 82.690 201.825 83.020 201.945 ;
        RECT 82.690 201.125 83.990 201.825 ;
        RECT 98.985 201.470 99.515 202.000 ;
        RECT 107.265 201.540 107.795 202.070 ;
        RECT 99.100 201.265 99.400 201.470 ;
        RECT 53.570 200.615 58.320 200.785 ;
        RECT 51.895 199.140 53.135 199.840 ;
        RECT 59.000 199.380 59.530 199.910 ;
        RECT 76.265 199.395 76.795 199.925 ;
        RECT 52.805 198.255 53.135 199.140 ;
        RECT 53.570 198.335 58.320 198.505 ;
        RECT 53.655 198.010 53.955 198.335 ;
        RECT 53.540 197.480 54.070 198.010 ;
        RECT 77.505 197.415 82.255 197.585 ;
        RECT 77.825 197.030 78.125 197.415 ;
        RECT 82.690 197.335 83.020 201.125 ;
        RECT 98.795 201.095 103.545 201.265 ;
        RECT 103.980 200.485 104.310 201.345 ;
        RECT 107.380 201.265 107.680 201.540 ;
        RECT 106.875 201.095 111.625 201.265 ;
        RECT 104.615 200.485 105.145 200.690 ;
        RECT 103.980 200.160 105.145 200.485 ;
        RECT 112.060 200.485 112.390 201.345 ;
        RECT 112.695 200.485 113.225 200.690 ;
        RECT 112.060 200.160 113.225 200.485 ;
        RECT 103.980 200.155 105.045 200.160 ;
        RECT 112.060 200.155 113.125 200.160 ;
        RECT 97.590 198.855 98.190 199.455 ;
        RECT 52.805 195.150 53.135 196.055 ;
        RECT 53.810 195.975 54.510 196.790 ;
        RECT 77.710 196.500 78.240 197.030 ;
        RECT 98.795 196.815 103.545 196.985 ;
        RECT 103.315 196.435 103.485 196.815 ;
        RECT 103.980 196.735 104.310 200.155 ;
        RECT 105.785 199.170 106.385 199.770 ;
        RECT 106.875 196.815 111.625 196.985 ;
        RECT 107.170 196.435 107.470 196.815 ;
        RECT 112.060 196.735 112.390 200.155 ;
        RECT 53.570 195.805 58.320 195.975 ;
        RECT 51.895 194.450 53.135 195.150 ;
        RECT 81.465 194.950 82.165 195.980 ;
        RECT 103.135 195.905 103.665 196.435 ;
        RECT 107.055 195.905 107.585 196.435 ;
        RECT 52.805 193.445 53.135 194.450 ;
        RECT 59.000 194.335 59.530 194.865 ;
        RECT 77.505 194.780 82.255 194.950 ;
        RECT 82.690 194.930 83.020 195.030 ;
        RECT 82.690 194.230 83.990 194.930 ;
        RECT 98.985 194.495 99.515 195.025 ;
        RECT 107.265 194.560 107.795 195.090 ;
        RECT 99.165 194.240 99.335 194.495 ;
        RECT 53.570 193.525 58.320 193.695 ;
        RECT 53.620 193.190 53.920 193.525 ;
        RECT 53.540 192.660 54.070 193.190 ;
        RECT 76.245 192.120 76.775 192.650 ;
        RECT 77.505 190.500 82.255 190.670 ;
        RECT 77.825 190.165 78.125 190.500 ;
        RECT 82.690 190.420 83.020 194.230 ;
        RECT 98.795 194.070 103.545 194.240 ;
        RECT 103.980 193.385 104.310 194.320 ;
        RECT 107.380 194.240 107.680 194.560 ;
        RECT 106.875 194.070 111.625 194.240 ;
        RECT 104.615 193.385 105.145 193.625 ;
        RECT 103.980 193.095 105.145 193.385 ;
        RECT 103.980 193.055 105.045 193.095 ;
        RECT 97.590 191.830 98.190 192.430 ;
        RECT 77.710 189.635 78.240 190.165 ;
        RECT 98.795 189.790 103.545 189.960 ;
        RECT 103.315 189.275 103.485 189.790 ;
        RECT 103.980 189.710 104.310 193.055 ;
        RECT 112.060 192.945 112.390 194.320 ;
        RECT 112.695 192.945 113.225 193.185 ;
        RECT 112.060 192.655 113.225 192.945 ;
        RECT 112.060 192.615 113.125 192.655 ;
        RECT 105.785 191.830 106.385 192.430 ;
        RECT 106.875 189.790 111.625 189.960 ;
        RECT 107.170 189.275 107.470 189.790 ;
        RECT 112.060 189.710 112.390 192.615 ;
        RECT 45.710 187.580 46.040 187.660 ;
        RECT 46.575 187.580 47.275 188.755 ;
        RECT 103.135 188.745 103.665 189.275 ;
        RECT 107.055 188.745 107.585 189.275 ;
        RECT 44.650 186.880 46.040 187.580 ;
        RECT 46.455 187.410 53.245 187.580 ;
        RECT 45.710 185.050 46.040 186.880 ;
        RECT 53.860 186.065 54.390 186.595 ;
        RECT 46.455 185.130 53.245 185.300 ;
        RECT 52.940 184.770 53.240 185.130 ;
        RECT 52.850 184.240 53.380 184.770 ;
        RECT 58.545 184.050 58.715 185.930 ;
        RECT 118.880 185.260 119.050 185.930 ;
        RECT 45.710 183.125 46.040 183.185 ;
        RECT 44.650 182.425 46.040 183.125 ;
        RECT 46.575 183.105 47.275 184.025 ;
        RECT 46.455 182.935 53.245 183.105 ;
        RECT 45.710 180.575 46.040 182.425 ;
        RECT 53.860 181.610 54.390 182.140 ;
        RECT 58.545 181.630 58.715 183.510 ;
        RECT 118.880 182.840 119.050 184.720 ;
        RECT 46.455 180.655 53.245 180.825 ;
        RECT 52.935 180.255 53.235 180.655 ;
        RECT 52.850 179.725 53.380 180.255 ;
        RECT 45.710 178.525 46.040 178.570 ;
        RECT 44.650 177.825 46.040 178.525 ;
        RECT 46.575 178.490 47.275 179.460 ;
        RECT 58.545 179.210 58.715 181.090 ;
        RECT 118.880 180.420 119.050 182.300 ;
        RECT 118.880 179.210 119.050 179.880 ;
        RECT 46.455 178.320 53.245 178.490 ;
        RECT 45.710 175.960 46.040 177.825 ;
        RECT 53.860 176.915 54.390 177.445 ;
        RECT 46.455 176.040 53.245 176.210 ;
        RECT 52.940 175.655 53.240 176.040 ;
        RECT 52.850 175.125 53.380 175.655 ;
        RECT 89.250 175.625 89.780 176.155 ;
        RECT 107.000 175.625 107.700 176.645 ;
        RECT 89.395 175.240 89.695 175.625 ;
        RECT 107.000 175.520 111.850 175.625 ;
        RECT 107.100 175.455 111.850 175.520 ;
        RECT 89.395 175.070 90.065 175.240 ;
        RECT 89.395 175.010 89.695 175.070 ;
        RECT 45.690 172.980 46.020 172.995 ;
        RECT 44.650 172.280 46.020 172.980 ;
        RECT 46.490 172.915 47.190 173.890 ;
        RECT 87.895 173.620 88.785 174.510 ;
        RECT 90.540 174.265 90.870 175.320 ;
        RECT 112.285 174.965 112.615 175.705 ;
        RECT 112.285 174.265 113.730 174.965 ;
        RECT 90.540 173.565 91.805 174.265 ;
        RECT 46.435 172.745 53.225 172.915 ;
        RECT 89.395 172.790 90.065 172.960 ;
        RECT 45.690 170.385 46.020 172.280 ;
        RECT 89.395 172.185 89.695 172.790 ;
        RECT 90.540 172.710 90.870 173.565 ;
        RECT 105.755 172.765 106.355 173.365 ;
        RECT 53.835 171.205 54.365 171.735 ;
        RECT 89.275 171.655 89.805 172.185 ;
        RECT 107.200 171.345 107.900 171.355 ;
        RECT 107.100 171.175 111.850 171.345 ;
        RECT 46.435 170.465 53.225 170.635 ;
        RECT 45.690 168.340 46.020 168.480 ;
        RECT 46.490 168.400 47.190 169.440 ;
        RECT 52.505 169.430 53.205 170.465 ;
        RECT 107.200 170.230 107.900 171.175 ;
        RECT 112.285 171.095 112.615 174.265 ;
        RECT 107.000 168.515 107.700 169.475 ;
        RECT 107.000 168.425 111.850 168.515 ;
        RECT 44.715 167.640 46.020 168.340 ;
        RECT 46.435 168.230 53.225 168.400 ;
        RECT 107.100 168.345 111.850 168.425 ;
        RECT 112.285 168.410 112.615 168.595 ;
        RECT 45.690 165.870 46.020 167.640 ;
        RECT 112.285 167.710 113.640 168.410 ;
        RECT 53.865 166.895 54.395 167.425 ;
        RECT 46.435 165.950 53.225 166.120 ;
        RECT 52.505 164.890 53.205 165.950 ;
        RECT 89.265 165.565 89.795 166.095 ;
        RECT 93.990 165.595 94.520 166.125 ;
        RECT 105.755 165.975 106.355 166.575 ;
        RECT 89.400 165.240 89.700 165.565 ;
        RECT 89.390 165.070 90.060 165.240 ;
        RECT 89.400 165.000 89.700 165.070 ;
        RECT 45.690 163.875 46.020 163.890 ;
        RECT 44.650 163.175 46.020 163.875 ;
        RECT 46.490 163.810 47.190 164.865 ;
        RECT 46.435 163.640 53.225 163.810 ;
        RECT 87.985 163.660 88.875 164.550 ;
        RECT 90.535 164.310 90.865 165.320 ;
        RECT 45.690 161.280 46.020 163.175 ;
        RECT 90.535 163.610 91.870 164.310 ;
        RECT 107.100 164.065 111.850 164.235 ;
        RECT 53.845 162.295 54.375 162.825 ;
        RECT 89.390 162.790 90.060 162.960 ;
        RECT 89.400 162.195 89.700 162.790 ;
        RECT 90.535 162.710 90.865 163.610 ;
        RECT 107.200 163.090 107.900 164.065 ;
        RECT 112.285 163.985 112.615 167.710 ;
        RECT 89.275 161.665 89.805 162.195 ;
        RECT 46.435 161.360 53.225 161.530 ;
        RECT 52.485 160.140 53.185 161.360 ;
        RECT 45.905 156.390 46.075 158.270 ;
        RECT 110.910 157.600 111.080 158.270 ;
        RECT 45.905 153.970 46.075 155.850 ;
        RECT 110.910 155.180 111.080 157.060 ;
        RECT 45.905 151.550 46.075 153.430 ;
        RECT 110.910 152.760 111.080 154.640 ;
        RECT 45.905 149.130 46.075 151.010 ;
        RECT 110.910 150.340 111.080 152.220 ;
        RECT 45.905 146.710 46.075 148.590 ;
        RECT 110.910 147.920 111.080 149.800 ;
        RECT 45.905 144.290 46.075 146.170 ;
        RECT 110.910 145.500 111.080 147.380 ;
        RECT 45.905 141.870 46.075 143.750 ;
        RECT 110.910 143.080 111.080 144.960 ;
        RECT 45.905 139.450 46.075 141.330 ;
        RECT 110.910 140.660 111.080 142.540 ;
        RECT 110.910 139.450 111.080 140.120 ;
        RECT 44.225 107.745 44.755 107.915 ;
        RECT 53.210 107.755 53.740 107.925 ;
        RECT 63.445 107.755 63.975 107.925 ;
        RECT 43.590 105.900 43.920 107.145 ;
        RECT 44.400 107.065 44.570 107.745 ;
        RECT 53.385 107.120 53.555 107.755 ;
        RECT 44.355 106.895 49.105 107.065 ;
        RECT 53.370 106.950 58.120 107.120 ;
        RECT 44.400 106.890 44.570 106.895 ;
        RECT 42.235 104.900 43.920 105.900 ;
        RECT 58.555 105.325 58.885 107.200 ;
        RECT 63.620 107.120 63.790 107.755 ;
        RECT 63.520 106.950 68.270 107.120 ;
        RECT 68.705 105.365 69.035 107.200 ;
        RECT 76.835 107.075 77.535 108.505 ;
        RECT 72.800 106.905 77.550 107.075 ;
        RECT 76.835 106.895 77.535 106.905 ;
        RECT 43.590 102.535 43.920 104.900 ;
        RECT 49.765 104.760 50.295 105.290 ;
        RECT 58.555 105.255 59.930 105.325 ;
        RECT 68.705 105.255 70.140 105.365 ;
        RECT 58.555 105.085 60.215 105.255 ;
        RECT 68.705 105.085 70.240 105.255 ;
        RECT 58.555 104.995 59.930 105.085 ;
        RECT 68.705 105.035 70.140 105.085 ;
        RECT 52.205 102.795 52.735 103.325 ;
        RECT 44.355 102.615 49.105 102.785 ;
        RECT 53.370 102.670 58.120 102.840 ;
        RECT 44.425 102.165 44.595 102.615 ;
        RECT 53.410 102.200 53.580 102.670 ;
        RECT 58.555 102.590 58.885 104.995 ;
        RECT 62.365 102.765 62.895 103.295 ;
        RECT 63.520 102.670 68.270 102.840 ;
        RECT 43.965 101.165 44.965 102.165 ;
        RECT 52.950 101.200 53.950 102.200 ;
        RECT 63.905 102.140 64.075 102.670 ;
        RECT 68.705 102.590 69.035 105.035 ;
        RECT 71.565 104.555 72.095 105.085 ;
        RECT 72.800 102.625 77.550 102.795 ;
        RECT 63.445 101.140 64.445 102.140 ;
        RECT 72.820 102.120 72.990 102.625 ;
        RECT 72.415 101.230 73.305 102.120 ;
        RECT 77.985 101.585 78.315 107.155 ;
        RECT 81.140 103.260 81.310 103.930 ;
        RECT 77.700 101.540 78.315 101.585 ;
        RECT 77.600 101.370 78.315 101.540 ;
        RECT 77.700 101.255 78.315 101.370 ;
        RECT 81.140 100.840 81.310 102.720 ;
        RECT 121.975 102.050 122.145 103.930 ;
        RECT 44.225 98.895 44.755 99.065 ;
        RECT 43.590 96.105 43.920 97.330 ;
        RECT 44.400 97.250 44.570 98.895 ;
        RECT 53.210 97.795 53.740 97.965 ;
        RECT 63.445 97.815 63.975 97.985 ;
        RECT 44.355 97.080 49.105 97.250 ;
        RECT 53.385 97.225 53.555 97.795 ;
        RECT 53.370 97.055 58.120 97.225 ;
        RECT 42.235 95.105 43.920 96.105 ;
        RECT 43.590 92.720 43.920 95.105 ;
        RECT 49.785 94.650 50.315 95.180 ;
        RECT 58.555 94.935 58.885 97.305 ;
        RECT 63.620 97.245 63.790 97.815 ;
        RECT 62.365 96.570 62.895 97.100 ;
        RECT 63.520 97.075 68.270 97.245 ;
        RECT 68.705 95.040 69.035 97.325 ;
        RECT 76.835 97.185 77.535 98.600 ;
        RECT 81.140 98.420 81.310 100.300 ;
        RECT 121.975 99.630 122.145 101.510 ;
        RECT 121.975 98.420 122.145 99.090 ;
        RECT 72.800 97.015 77.550 97.185 ;
        RECT 76.835 96.990 77.535 97.015 ;
        RECT 58.555 94.905 59.975 94.935 ;
        RECT 68.705 94.905 70.140 95.040 ;
        RECT 58.555 94.735 60.215 94.905 ;
        RECT 68.705 94.735 70.240 94.905 ;
        RECT 58.555 94.605 59.975 94.735 ;
        RECT 68.705 94.710 70.140 94.735 ;
        RECT 44.355 92.800 49.105 92.970 ;
        RECT 52.205 92.865 52.735 93.395 ;
        RECT 44.425 92.255 44.595 92.800 ;
        RECT 53.370 92.775 58.120 92.945 ;
        RECT 53.410 92.290 53.580 92.775 ;
        RECT 58.555 92.695 58.885 94.605 ;
        RECT 63.520 92.795 68.270 92.965 ;
        RECT 43.965 91.255 44.965 92.255 ;
        RECT 52.950 91.290 53.950 92.290 ;
        RECT 63.905 92.245 64.075 92.795 ;
        RECT 68.705 92.715 69.035 94.710 ;
        RECT 71.585 94.590 72.115 95.120 ;
        RECT 72.800 92.735 77.550 92.905 ;
        RECT 63.445 91.245 64.445 92.245 ;
        RECT 72.820 92.220 72.990 92.735 ;
        RECT 72.415 91.330 73.305 92.220 ;
        RECT 77.985 92.070 78.315 97.265 ;
        RECT 91.430 94.530 91.960 95.060 ;
        RECT 94.635 94.465 95.635 95.465 ;
        RECT 110.465 95.125 110.995 95.655 ;
        RECT 96.325 94.685 96.855 94.855 ;
        RECT 92.730 92.765 93.730 93.740 ;
        RECT 94.395 93.580 94.925 93.605 ;
        RECT 94.395 93.435 95.010 93.580 ;
        RECT 94.765 93.410 95.010 93.435 ;
        RECT 92.730 92.740 94.570 92.765 ;
        RECT 93.305 92.595 94.570 92.740 ;
        RECT 77.700 92.020 78.315 92.070 ;
        RECT 77.600 91.850 78.315 92.020 ;
        RECT 77.700 91.740 78.315 91.850 ;
        RECT 91.700 91.175 92.700 92.175 ;
        RECT 94.400 92.105 94.570 92.595 ;
        RECT 94.840 92.520 95.010 93.410 ;
        RECT 95.360 93.140 95.530 94.465 ;
        RECT 96.505 93.780 96.675 94.685 ;
        RECT 112.965 94.465 113.965 95.465 ;
        RECT 114.655 94.685 115.185 94.855 ;
        RECT 96.200 93.610 100.950 93.780 ;
        RECT 96.200 93.140 100.950 93.150 ;
        RECT 95.360 92.980 100.950 93.140 ;
        RECT 95.360 92.970 96.330 92.980 ;
        RECT 101.385 92.615 101.715 93.860 ;
        RECT 102.765 92.615 103.765 93.055 ;
        RECT 111.060 92.765 112.060 93.740 ;
        RECT 112.725 93.580 113.255 93.605 ;
        RECT 112.725 93.435 113.340 93.580 ;
        RECT 113.095 93.410 113.340 93.435 ;
        RECT 111.060 92.740 112.900 92.765 ;
        RECT 94.840 92.350 100.950 92.520 ;
        RECT 101.385 92.285 103.765 92.615 ;
        RECT 111.635 92.595 112.900 92.740 ;
        RECT 94.400 91.935 95.900 92.105 ;
        RECT 93.345 91.765 93.960 91.935 ;
        RECT 93.790 91.700 93.960 91.765 ;
        RECT 95.730 91.890 95.900 91.935 ;
        RECT 95.730 91.720 100.950 91.890 ;
        RECT 93.790 91.530 95.440 91.700 ;
        RECT 95.270 91.460 95.440 91.530 ;
        RECT 95.270 91.290 95.915 91.460 ;
        RECT 92.530 91.070 92.700 91.175 ;
        RECT 95.745 91.260 95.915 91.290 ;
        RECT 95.745 91.090 100.950 91.260 ;
        RECT 92.530 90.900 95.335 91.070 ;
        RECT 89.350 89.670 90.350 90.670 ;
        RECT 95.165 90.630 95.335 90.900 ;
        RECT 91.590 90.420 94.975 90.590 ;
        RECT 95.165 90.460 100.950 90.630 ;
        RECT 91.590 90.355 91.760 90.420 ;
        RECT 91.230 90.185 91.760 90.355 ;
        RECT 92.385 89.895 94.250 90.065 ;
        RECT 88.030 89.455 88.560 89.540 ;
        RECT 88.030 89.285 88.820 89.455 ;
        RECT 88.650 88.885 88.820 89.285 ;
        RECT 90.000 89.345 90.170 89.670 ;
        RECT 92.385 89.345 92.555 89.895 ;
        RECT 90.000 89.175 92.555 89.345 ;
        RECT 94.080 89.370 94.250 89.895 ;
        RECT 94.805 90.000 94.975 90.420 ;
        RECT 94.805 89.830 100.950 90.000 ;
        RECT 94.080 89.200 100.950 89.370 ;
        RECT 89.640 88.885 91.915 88.910 ;
        RECT 53.210 88.025 53.740 88.195 ;
        RECT 63.445 88.150 63.975 88.320 ;
        RECT 44.225 87.675 44.755 87.845 ;
        RECT 43.590 86.745 43.920 87.170 ;
        RECT 44.400 87.090 44.570 87.675 ;
        RECT 53.395 87.180 53.565 88.025 ;
        RECT 63.630 87.305 63.800 88.150 ;
        RECT 44.355 86.920 49.105 87.090 ;
        RECT 53.370 87.010 58.120 87.180 ;
        RECT 42.235 85.745 43.920 86.745 ;
        RECT 43.590 82.560 43.920 85.745 ;
        RECT 49.765 84.575 50.295 85.105 ;
        RECT 58.555 84.950 58.885 87.260 ;
        RECT 63.520 87.135 68.270 87.305 ;
        RECT 62.365 86.565 62.895 87.095 ;
        RECT 68.705 85.100 69.035 87.385 ;
        RECT 76.785 87.350 77.485 88.790 ;
        RECT 88.650 88.740 91.915 88.885 ;
        RECT 88.650 88.715 89.810 88.740 ;
        RECT 91.745 88.570 100.950 88.740 ;
        RECT 86.135 88.110 87.135 88.510 ;
        RECT 86.135 87.940 100.950 88.110 ;
        RECT 86.135 87.510 87.135 87.940 ;
        RECT 96.200 87.450 100.950 87.480 ;
        RECT 72.755 87.180 77.505 87.350 ;
        RECT 68.705 85.045 70.140 85.100 ;
        RECT 58.555 84.885 60.020 84.950 ;
        RECT 58.555 84.715 60.215 84.885 ;
        RECT 68.705 84.875 70.240 85.045 ;
        RECT 68.705 84.770 70.140 84.875 ;
        RECT 71.525 84.830 72.055 85.360 ;
        RECT 58.555 84.620 60.020 84.715 ;
        RECT 52.205 82.815 52.735 83.345 ;
        RECT 44.355 82.640 49.105 82.810 ;
        RECT 53.370 82.730 58.120 82.900 ;
        RECT 44.425 82.100 44.595 82.640 ;
        RECT 53.410 82.275 53.580 82.730 ;
        RECT 58.555 82.650 58.885 84.620 ;
        RECT 63.520 82.855 68.270 83.025 ;
        RECT 63.905 82.390 64.075 82.855 ;
        RECT 68.705 82.775 69.035 84.770 ;
        RECT 72.755 82.900 77.505 83.070 ;
        RECT 72.760 82.540 72.930 82.900 ;
        RECT 43.965 81.100 44.965 82.100 ;
        RECT 52.950 81.275 53.950 82.275 ;
        RECT 63.445 81.390 64.445 82.390 ;
        RECT 72.490 81.540 73.490 82.540 ;
        RECT 77.940 81.665 78.270 87.430 ;
        RECT 94.660 87.310 100.950 87.450 ;
        RECT 94.660 87.280 96.415 87.310 ;
        RECT 94.660 87.180 94.830 87.280 ;
        RECT 88.030 87.010 94.830 87.180 ;
        RECT 95.225 86.850 96.365 86.865 ;
        RECT 95.225 86.695 100.950 86.850 ;
        RECT 95.225 86.645 95.395 86.695 ;
        RECT 96.200 86.680 100.950 86.695 ;
        RECT 89.085 86.475 95.395 86.645 ;
        RECT 89.085 86.130 89.255 86.475 ;
        RECT 96.200 86.200 100.950 86.220 ;
        RECT 95.685 86.160 100.950 86.200 ;
        RECT 88.670 85.130 89.670 86.130 ;
        RECT 90.810 86.050 100.950 86.160 ;
        RECT 90.810 86.030 96.355 86.050 ;
        RECT 90.810 85.990 95.855 86.030 ;
        RECT 90.810 85.715 90.980 85.990 ;
        RECT 90.365 85.545 90.980 85.715 ;
        RECT 91.465 85.420 100.950 85.590 ;
        RECT 91.465 84.705 91.635 85.420 ;
        RECT 92.930 84.790 100.950 84.960 ;
        RECT 90.745 83.705 91.745 84.705 ;
        RECT 92.930 84.195 93.100 84.790 ;
        RECT 92.470 84.025 93.100 84.195 ;
        RECT 92.650 83.985 93.100 84.025 ;
        RECT 93.640 84.160 100.950 84.330 ;
        RECT 93.640 83.290 93.810 84.160 ;
        RECT 91.620 83.120 93.810 83.290 ;
        RECT 94.250 83.530 100.950 83.700 ;
        RECT 91.620 82.760 91.790 83.120 ;
        RECT 90.745 82.175 91.790 82.760 ;
        RECT 94.250 82.440 94.420 83.530 ;
        RECT 92.855 82.370 94.420 82.440 ;
        RECT 92.675 82.270 94.420 82.370 ;
        RECT 94.870 82.900 100.950 83.070 ;
        RECT 92.675 82.200 93.205 82.270 ;
        RECT 90.745 81.760 91.745 82.175 ;
        RECT 94.870 81.885 95.040 82.900 ;
        RECT 77.565 81.500 78.270 81.665 ;
        RECT 93.810 81.715 95.040 81.885 ;
        RECT 95.360 82.270 100.950 82.440 ;
        RECT 77.565 81.495 78.095 81.500 ;
        RECT 93.810 81.220 93.980 81.715 ;
        RECT 93.015 80.220 94.015 81.220 ;
        RECT 95.360 80.945 95.530 82.270 ;
        RECT 96.200 81.640 100.950 81.810 ;
        RECT 96.585 81.220 96.755 81.640 ;
        RECT 101.385 81.560 101.715 92.285 ;
        RECT 102.765 92.055 103.765 92.285 ;
        RECT 110.030 91.175 111.030 92.175 ;
        RECT 112.730 92.105 112.900 92.595 ;
        RECT 113.170 92.520 113.340 93.410 ;
        RECT 113.690 93.140 113.860 94.465 ;
        RECT 114.835 93.780 115.005 94.685 ;
        RECT 114.545 93.610 119.295 93.780 ;
        RECT 114.545 93.140 119.295 93.150 ;
        RECT 113.690 92.980 119.295 93.140 ;
        RECT 113.690 92.970 114.660 92.980 ;
        RECT 113.170 92.350 119.295 92.520 ;
        RECT 112.730 91.935 114.230 92.105 ;
        RECT 111.675 91.765 112.290 91.935 ;
        RECT 112.120 91.700 112.290 91.765 ;
        RECT 114.060 91.890 114.230 91.935 ;
        RECT 114.060 91.720 119.295 91.890 ;
        RECT 112.120 91.530 113.770 91.700 ;
        RECT 113.600 91.460 113.770 91.530 ;
        RECT 113.600 91.290 114.245 91.460 ;
        RECT 110.860 91.070 111.030 91.175 ;
        RECT 114.075 91.260 114.245 91.290 ;
        RECT 114.075 91.090 119.295 91.260 ;
        RECT 110.860 90.900 113.665 91.070 ;
        RECT 107.680 89.670 108.680 90.670 ;
        RECT 113.495 90.630 113.665 90.900 ;
        RECT 109.920 90.420 113.305 90.590 ;
        RECT 113.495 90.460 119.295 90.630 ;
        RECT 109.920 90.355 110.090 90.420 ;
        RECT 109.560 90.185 110.090 90.355 ;
        RECT 110.715 89.895 112.580 90.065 ;
        RECT 106.360 89.455 106.890 89.540 ;
        RECT 106.360 89.285 107.150 89.455 ;
        RECT 106.980 88.885 107.150 89.285 ;
        RECT 108.330 89.345 108.500 89.670 ;
        RECT 110.715 89.345 110.885 89.895 ;
        RECT 108.330 89.175 110.885 89.345 ;
        RECT 112.410 89.370 112.580 89.895 ;
        RECT 113.135 90.000 113.305 90.420 ;
        RECT 113.135 89.830 119.295 90.000 ;
        RECT 112.410 89.200 119.295 89.370 ;
        RECT 107.970 88.885 110.245 88.910 ;
        RECT 106.980 88.740 110.245 88.885 ;
        RECT 106.980 88.715 108.140 88.740 ;
        RECT 110.075 88.570 119.295 88.740 ;
        RECT 104.465 88.110 105.465 88.530 ;
        RECT 119.730 88.485 120.060 93.860 ;
        RECT 104.465 87.940 119.295 88.110 ;
        RECT 104.465 87.530 105.465 87.940 ;
        RECT 119.730 87.785 121.175 88.485 ;
        RECT 114.545 87.450 119.295 87.480 ;
        RECT 112.990 87.310 119.295 87.450 ;
        RECT 112.990 87.280 114.745 87.310 ;
        RECT 112.990 87.180 113.160 87.280 ;
        RECT 106.360 87.010 113.160 87.180 ;
        RECT 113.555 86.850 114.695 86.865 ;
        RECT 113.555 86.695 119.295 86.850 ;
        RECT 113.555 86.645 113.725 86.695 ;
        RECT 114.545 86.680 119.295 86.695 ;
        RECT 107.415 86.475 113.725 86.645 ;
        RECT 107.415 86.130 107.585 86.475 ;
        RECT 114.545 86.200 119.295 86.220 ;
        RECT 114.015 86.160 119.295 86.200 ;
        RECT 107.000 85.130 108.000 86.130 ;
        RECT 109.140 86.050 119.295 86.160 ;
        RECT 109.140 86.030 114.685 86.050 ;
        RECT 109.140 85.990 114.185 86.030 ;
        RECT 109.140 85.715 109.310 85.990 ;
        RECT 108.695 85.545 109.310 85.715 ;
        RECT 109.795 85.420 119.295 85.590 ;
        RECT 109.795 84.705 109.965 85.420 ;
        RECT 111.260 84.790 119.295 84.960 ;
        RECT 109.075 83.705 110.075 84.705 ;
        RECT 111.260 84.195 111.430 84.790 ;
        RECT 110.800 84.025 111.430 84.195 ;
        RECT 110.980 83.985 111.430 84.025 ;
        RECT 111.970 84.160 119.295 84.330 ;
        RECT 111.970 83.290 112.140 84.160 ;
        RECT 109.950 83.120 112.140 83.290 ;
        RECT 112.580 83.530 119.295 83.700 ;
        RECT 109.950 82.760 110.120 83.120 ;
        RECT 109.075 82.175 110.120 82.760 ;
        RECT 112.580 82.440 112.750 83.530 ;
        RECT 111.185 82.370 112.750 82.440 ;
        RECT 111.005 82.270 112.750 82.370 ;
        RECT 113.200 82.900 119.295 83.070 ;
        RECT 111.005 82.200 111.535 82.270 ;
        RECT 109.075 81.760 110.075 82.175 ;
        RECT 113.200 81.885 113.370 82.900 ;
        RECT 112.140 81.715 113.370 81.885 ;
        RECT 113.690 82.270 119.295 82.440 ;
        RECT 112.140 81.220 112.310 81.715 ;
        RECT 94.935 80.910 95.530 80.945 ;
        RECT 94.755 80.775 95.530 80.910 ;
        RECT 94.755 80.740 95.285 80.775 ;
        RECT 96.170 80.220 97.170 81.220 ;
        RECT 111.345 80.220 112.345 81.220 ;
        RECT 113.690 80.945 113.860 82.270 ;
        RECT 114.545 81.640 119.295 81.810 ;
        RECT 114.915 81.220 115.085 81.640 ;
        RECT 119.730 81.560 120.060 87.785 ;
        RECT 113.265 80.910 113.860 80.945 ;
        RECT 113.085 80.775 113.860 80.910 ;
        RECT 113.085 80.740 113.615 80.775 ;
        RECT 114.500 80.220 115.500 81.220 ;
        RECT 44.225 78.600 44.755 78.770 ;
        RECT 43.590 76.175 43.920 78.105 ;
        RECT 44.400 78.025 44.570 78.600 ;
        RECT 53.210 78.590 53.740 78.760 ;
        RECT 63.445 78.635 63.975 78.805 ;
        RECT 44.355 77.855 49.105 78.025 ;
        RECT 53.385 77.980 53.555 78.590 ;
        RECT 52.205 77.395 52.735 77.925 ;
        RECT 53.370 77.810 58.120 77.980 ;
        RECT 41.865 75.175 43.920 76.175 ;
        RECT 58.555 76.000 58.885 78.060 ;
        RECT 63.620 77.885 63.790 78.635 ;
        RECT 77.035 78.490 77.565 78.495 ;
        RECT 76.855 78.325 77.565 78.490 ;
        RECT 62.365 77.300 62.895 77.830 ;
        RECT 63.520 77.715 68.270 77.885 ;
        RECT 58.555 75.950 59.985 76.000 ;
        RECT 49.785 75.375 50.315 75.905 ;
        RECT 58.555 75.780 60.215 75.950 ;
        RECT 58.555 75.670 59.985 75.780 ;
        RECT 68.705 75.770 69.035 77.965 ;
        RECT 76.855 77.790 77.555 78.325 ;
        RECT 72.800 77.620 77.555 77.790 ;
        RECT 76.855 77.605 77.555 77.620 ;
        RECT 68.705 75.720 69.915 75.770 ;
        RECT 43.590 73.495 43.920 75.175 ;
        RECT 44.355 73.575 49.105 73.745 ;
        RECT 44.425 73.095 44.595 73.575 ;
        RECT 53.370 73.530 58.120 73.700 ;
        RECT 43.965 72.095 44.965 73.095 ;
        RECT 53.410 73.070 53.580 73.530 ;
        RECT 58.555 73.450 58.885 75.670 ;
        RECT 68.705 75.550 70.240 75.720 ;
        RECT 68.705 75.440 69.915 75.550 ;
        RECT 63.520 73.435 68.270 73.605 ;
        RECT 63.905 73.215 64.075 73.435 ;
        RECT 68.705 73.355 69.035 75.440 ;
        RECT 71.545 75.130 72.075 75.660 ;
        RECT 72.810 73.510 72.980 73.530 ;
        RECT 72.800 73.340 77.550 73.510 ;
        RECT 52.950 72.070 53.950 73.070 ;
        RECT 63.445 72.215 64.445 73.215 ;
        RECT 72.810 72.915 72.980 73.340 ;
        RECT 72.085 71.915 73.085 72.915 ;
        RECT 77.985 72.225 78.315 77.870 ;
        RECT 91.120 76.145 91.650 76.675 ;
        RECT 94.395 76.175 95.395 77.175 ;
        RECT 96.035 76.395 96.565 76.565 ;
        RECT 92.440 74.475 93.440 75.450 ;
        RECT 94.105 75.290 94.635 75.315 ;
        RECT 94.105 75.145 94.720 75.290 ;
        RECT 94.475 75.120 94.720 75.145 ;
        RECT 92.440 74.450 94.280 74.475 ;
        RECT 93.015 74.305 94.280 74.450 ;
        RECT 91.410 72.885 92.410 73.885 ;
        RECT 94.110 73.815 94.280 74.305 ;
        RECT 94.550 74.230 94.720 75.120 ;
        RECT 95.070 74.850 95.240 76.175 ;
        RECT 96.215 75.490 96.385 76.395 ;
        RECT 109.770 75.770 110.300 76.300 ;
        RECT 112.995 75.930 113.995 76.930 ;
        RECT 114.685 76.150 115.215 76.320 ;
        RECT 95.895 75.320 100.645 75.490 ;
        RECT 95.895 74.850 100.645 74.860 ;
        RECT 95.070 74.690 100.645 74.850 ;
        RECT 95.070 74.680 96.040 74.690 ;
        RECT 94.550 74.060 100.645 74.230 ;
        RECT 94.110 73.645 95.610 73.815 ;
        RECT 93.055 73.475 93.670 73.645 ;
        RECT 93.500 73.410 93.670 73.475 ;
        RECT 95.440 73.600 95.610 73.645 ;
        RECT 95.440 73.430 100.645 73.600 ;
        RECT 93.500 73.240 95.150 73.410 ;
        RECT 94.980 73.170 95.150 73.240 ;
        RECT 94.980 73.000 95.625 73.170 ;
        RECT 92.240 72.780 92.410 72.885 ;
        RECT 95.455 72.970 95.625 73.000 ;
        RECT 95.455 72.800 100.645 72.970 ;
        RECT 92.240 72.610 95.045 72.780 ;
        RECT 77.695 71.895 78.315 72.225 ;
        RECT 89.060 71.380 90.060 72.380 ;
        RECT 94.875 72.340 95.045 72.610 ;
        RECT 91.300 72.130 94.685 72.300 ;
        RECT 94.875 72.170 100.645 72.340 ;
        RECT 91.300 72.065 91.470 72.130 ;
        RECT 90.940 71.895 91.470 72.065 ;
        RECT 92.095 71.605 93.960 71.775 ;
        RECT 87.740 71.165 88.270 71.250 ;
        RECT 87.740 70.995 88.530 71.165 ;
        RECT 49.275 70.765 50.340 70.860 ;
        RECT 49.275 70.595 50.440 70.765 ;
        RECT 88.360 70.595 88.530 70.995 ;
        RECT 89.710 71.055 89.880 71.380 ;
        RECT 92.095 71.055 92.265 71.605 ;
        RECT 89.710 70.885 92.265 71.055 ;
        RECT 93.790 71.080 93.960 71.605 ;
        RECT 94.515 71.710 94.685 72.130 ;
        RECT 94.515 71.540 100.645 71.710 ;
        RECT 93.790 70.910 100.645 71.080 ;
        RECT 89.350 70.595 91.625 70.620 ;
        RECT 49.275 70.530 50.340 70.595 ;
        RECT 49.275 66.280 49.605 70.530 ;
        RECT 50.040 69.810 50.210 70.530 ;
        RECT 88.360 70.450 91.625 70.595 ;
        RECT 88.360 70.425 89.520 70.450 ;
        RECT 91.455 70.280 100.645 70.450 ;
        RECT 85.845 69.820 86.845 70.240 ;
        RECT 50.030 69.640 55.800 69.810 ;
        RECT 85.845 69.650 100.645 69.820 ;
        RECT 85.845 69.240 86.845 69.650 ;
        RECT 95.895 69.160 100.645 69.190 ;
        RECT 94.370 69.020 100.645 69.160 ;
        RECT 94.370 68.990 96.125 69.020 ;
        RECT 94.370 68.890 94.540 68.990 ;
        RECT 87.740 68.720 94.540 68.890 ;
        RECT 94.935 68.560 96.075 68.575 ;
        RECT 73.830 68.265 74.360 68.440 ;
        RECT 94.935 68.405 100.645 68.560 ;
        RECT 94.935 68.355 95.105 68.405 ;
        RECT 95.895 68.390 100.645 68.405 ;
        RECT 73.830 68.095 81.840 68.265 ;
        RECT 73.830 67.910 74.360 68.095 ;
        RECT 62.085 67.795 62.815 67.800 ;
        RECT 61.905 67.785 62.815 67.795 ;
        RECT 56.440 67.120 56.970 67.650 ;
        RECT 61.905 67.630 69.485 67.785 ;
        RECT 61.905 67.625 62.435 67.630 ;
        RECT 62.695 67.615 69.485 67.630 ;
        RECT 59.755 66.705 69.485 66.875 ;
        RECT 50.030 66.510 55.800 66.530 ;
        RECT 50.020 66.360 55.800 66.510 ;
        RECT 50.020 65.895 50.190 66.360 ;
        RECT 49.560 64.895 50.560 65.895 ;
        RECT 59.755 65.055 59.925 66.705 ;
        RECT 62.085 65.975 62.945 65.980 ;
        RECT 61.905 65.965 62.945 65.975 ;
        RECT 61.905 65.810 69.485 65.965 ;
        RECT 61.905 65.805 62.435 65.810 ;
        RECT 62.695 65.795 69.485 65.810 ;
        RECT 59.755 64.885 69.485 65.055 ;
        RECT 49.275 64.225 50.340 64.255 ;
        RECT 49.275 64.055 50.440 64.225 ;
        RECT 49.275 63.925 50.340 64.055 ;
        RECT 49.275 59.590 49.605 63.925 ;
        RECT 50.030 63.120 50.200 63.925 ;
        RECT 59.755 63.235 59.925 64.885 ;
        RECT 62.085 64.155 62.925 64.160 ;
        RECT 61.905 64.145 62.925 64.155 ;
        RECT 61.905 63.990 69.485 64.145 ;
        RECT 61.905 63.985 62.435 63.990 ;
        RECT 62.695 63.975 69.485 63.990 ;
        RECT 50.030 62.950 55.800 63.120 ;
        RECT 59.755 63.065 69.485 63.235 ;
        RECT 56.460 61.785 56.990 62.315 ;
        RECT 59.755 61.415 59.925 63.065 ;
        RECT 61.915 62.325 62.815 62.340 ;
        RECT 61.915 62.170 69.485 62.325 ;
        RECT 62.695 62.155 69.485 62.170 ;
        RECT 59.755 61.245 69.485 61.415 ;
        RECT 50.030 59.820 55.800 59.840 ;
        RECT 50.020 59.670 55.800 59.820 ;
        RECT 50.020 59.205 50.190 59.670 ;
        RECT 59.755 59.595 59.925 61.245 ;
        RECT 61.915 60.505 62.445 60.515 ;
        RECT 61.915 60.345 69.485 60.505 ;
        RECT 62.095 60.335 69.485 60.345 ;
        RECT 59.755 59.425 69.485 59.595 ;
        RECT 49.560 58.205 50.560 59.205 ;
        RECT 59.755 57.775 59.925 59.425 ;
        RECT 62.095 58.690 62.960 58.700 ;
        RECT 61.915 58.685 62.960 58.690 ;
        RECT 61.915 58.530 69.485 58.685 ;
        RECT 61.915 58.520 62.445 58.530 ;
        RECT 62.695 58.515 69.485 58.530 ;
        RECT 59.755 57.605 69.485 57.775 ;
        RECT 49.275 57.530 50.340 57.600 ;
        RECT 49.275 57.360 50.440 57.530 ;
        RECT 49.275 57.270 50.340 57.360 ;
        RECT 49.275 52.900 49.605 57.270 ;
        RECT 50.035 56.430 50.205 57.270 ;
        RECT 59.755 56.765 59.925 57.605 ;
        RECT 61.905 56.865 62.950 56.880 ;
        RECT 60.325 56.765 60.595 56.850 ;
        RECT 59.755 56.595 60.595 56.765 ;
        RECT 61.905 56.710 69.485 56.865 ;
        RECT 62.695 56.695 69.485 56.710 ;
        RECT 50.030 56.260 55.800 56.430 ;
        RECT 59.755 55.955 59.925 56.595 ;
        RECT 60.325 56.520 60.595 56.595 ;
        RECT 59.755 55.785 69.485 55.955 ;
        RECT 59.755 55.055 59.925 55.785 ;
        RECT 62.180 55.060 62.375 55.175 ;
        RECT 62.180 55.055 62.910 55.060 ;
        RECT 59.610 54.885 60.140 55.055 ;
        RECT 61.915 55.045 62.910 55.055 ;
        RECT 61.915 54.890 69.485 55.045 ;
        RECT 69.900 55.030 70.230 67.865 ;
        RECT 72.630 66.815 81.840 66.985 ;
        RECT 72.680 64.425 72.850 66.815 ;
        RECT 73.830 65.705 74.360 65.925 ;
        RECT 73.830 65.535 81.840 65.705 ;
        RECT 73.830 65.395 74.360 65.535 ;
        RECT 72.680 64.255 81.840 64.425 ;
        RECT 72.680 61.865 72.850 64.255 ;
        RECT 73.830 63.145 74.360 63.320 ;
        RECT 73.830 62.975 81.840 63.145 ;
        RECT 73.830 62.790 74.360 62.975 ;
        RECT 72.680 61.695 81.840 61.865 ;
        RECT 72.680 59.305 72.850 61.695 ;
        RECT 73.830 60.585 74.360 60.790 ;
        RECT 73.830 60.415 81.840 60.585 ;
        RECT 73.830 60.260 74.360 60.415 ;
        RECT 72.680 59.135 81.840 59.305 ;
        RECT 72.680 56.745 72.850 59.135 ;
        RECT 73.830 58.025 74.360 58.145 ;
        RECT 73.830 57.855 81.840 58.025 ;
        RECT 73.830 57.615 74.360 57.855 ;
        RECT 72.680 56.575 81.840 56.745 ;
        RECT 72.680 56.165 72.850 56.575 ;
        RECT 72.680 56.015 72.955 56.165 ;
        RECT 72.685 55.835 72.955 56.015 ;
        RECT 61.915 54.885 62.445 54.890 ;
        RECT 62.695 54.875 69.485 54.890 ;
        RECT 69.880 54.795 70.230 55.030 ;
        RECT 72.710 55.000 72.880 55.835 ;
        RECT 73.830 55.465 74.360 55.670 ;
        RECT 73.830 55.295 81.840 55.465 ;
        RECT 73.830 55.140 74.360 55.295 ;
        RECT 82.255 55.215 82.585 68.345 ;
        RECT 88.795 68.185 95.105 68.355 ;
        RECT 88.795 67.840 88.965 68.185 ;
        RECT 95.895 67.910 100.645 67.930 ;
        RECT 95.395 67.870 100.645 67.910 ;
        RECT 88.380 66.840 89.380 67.840 ;
        RECT 90.520 67.760 100.645 67.870 ;
        RECT 90.520 67.740 96.065 67.760 ;
        RECT 90.520 67.700 95.565 67.740 ;
        RECT 90.520 67.425 90.690 67.700 ;
        RECT 90.075 67.255 90.690 67.425 ;
        RECT 91.175 67.130 100.645 67.300 ;
        RECT 91.175 66.415 91.345 67.130 ;
        RECT 92.640 66.500 100.645 66.670 ;
        RECT 90.455 65.415 91.455 66.415 ;
        RECT 92.640 65.905 92.810 66.500 ;
        RECT 92.180 65.735 92.810 65.905 ;
        RECT 92.360 65.695 92.810 65.735 ;
        RECT 93.350 65.870 100.645 66.040 ;
        RECT 93.350 65.000 93.520 65.870 ;
        RECT 91.330 64.830 93.520 65.000 ;
        RECT 93.960 65.240 100.645 65.410 ;
        RECT 91.330 64.470 91.500 64.830 ;
        RECT 90.455 63.885 91.500 64.470 ;
        RECT 93.960 64.150 94.130 65.240 ;
        RECT 92.565 64.080 94.130 64.150 ;
        RECT 92.385 63.980 94.130 64.080 ;
        RECT 94.580 64.610 100.645 64.780 ;
        RECT 92.385 63.910 92.915 63.980 ;
        RECT 90.455 63.470 91.455 63.885 ;
        RECT 94.580 63.595 94.750 64.610 ;
        RECT 101.080 64.325 101.410 75.570 ;
        RECT 111.090 74.230 112.090 75.205 ;
        RECT 112.755 75.045 113.285 75.070 ;
        RECT 112.755 74.900 113.370 75.045 ;
        RECT 113.125 74.875 113.370 74.900 ;
        RECT 111.090 74.205 112.930 74.230 ;
        RECT 111.665 74.060 112.930 74.205 ;
        RECT 110.060 72.640 111.060 73.640 ;
        RECT 112.760 73.570 112.930 74.060 ;
        RECT 113.200 73.985 113.370 74.875 ;
        RECT 113.720 74.605 113.890 75.930 ;
        RECT 114.865 75.245 115.035 76.150 ;
        RECT 114.550 75.075 119.300 75.245 ;
        RECT 114.550 74.605 119.300 74.615 ;
        RECT 113.720 74.445 119.300 74.605 ;
        RECT 113.720 74.435 114.690 74.445 ;
        RECT 113.200 73.815 119.300 73.985 ;
        RECT 112.760 73.400 114.260 73.570 ;
        RECT 111.705 73.230 112.320 73.400 ;
        RECT 112.150 73.165 112.320 73.230 ;
        RECT 114.090 73.355 114.260 73.400 ;
        RECT 114.090 73.185 119.300 73.355 ;
        RECT 112.150 72.995 113.800 73.165 ;
        RECT 113.630 72.925 113.800 72.995 ;
        RECT 113.630 72.755 114.275 72.925 ;
        RECT 110.890 72.535 111.060 72.640 ;
        RECT 114.105 72.725 114.275 72.755 ;
        RECT 114.105 72.555 119.300 72.725 ;
        RECT 110.890 72.365 113.695 72.535 ;
        RECT 107.710 71.135 108.710 72.135 ;
        RECT 113.525 72.095 113.695 72.365 ;
        RECT 109.950 71.885 113.335 72.055 ;
        RECT 113.525 71.925 119.300 72.095 ;
        RECT 109.950 71.820 110.120 71.885 ;
        RECT 109.590 71.650 110.120 71.820 ;
        RECT 110.745 71.360 112.610 71.530 ;
        RECT 106.390 70.920 106.920 71.005 ;
        RECT 106.390 70.750 107.180 70.920 ;
        RECT 107.010 70.350 107.180 70.750 ;
        RECT 108.360 70.810 108.530 71.135 ;
        RECT 110.745 70.810 110.915 71.360 ;
        RECT 108.360 70.640 110.915 70.810 ;
        RECT 112.440 70.835 112.610 71.360 ;
        RECT 113.165 71.465 113.335 71.885 ;
        RECT 113.165 71.295 119.300 71.465 ;
        RECT 112.440 70.665 119.300 70.835 ;
        RECT 108.000 70.350 110.275 70.375 ;
        RECT 107.010 70.205 110.275 70.350 ;
        RECT 107.010 70.180 108.170 70.205 ;
        RECT 110.105 70.035 119.300 70.205 ;
        RECT 104.495 69.575 105.495 70.010 ;
        RECT 119.735 69.880 120.065 75.325 ;
        RECT 104.495 69.405 119.300 69.575 ;
        RECT 104.495 69.010 105.495 69.405 ;
        RECT 119.735 69.180 120.900 69.880 ;
        RECT 114.550 68.915 119.300 68.945 ;
        RECT 113.020 68.775 119.300 68.915 ;
        RECT 113.020 68.745 114.775 68.775 ;
        RECT 113.020 68.645 113.190 68.745 ;
        RECT 106.390 68.475 113.190 68.645 ;
        RECT 113.585 68.315 114.725 68.330 ;
        RECT 113.585 68.160 119.300 68.315 ;
        RECT 113.585 68.110 113.755 68.160 ;
        RECT 114.550 68.145 119.300 68.160 ;
        RECT 107.445 67.940 113.755 68.110 ;
        RECT 107.445 67.595 107.615 67.940 ;
        RECT 114.550 67.665 119.300 67.685 ;
        RECT 114.045 67.625 119.300 67.665 ;
        RECT 107.030 66.595 108.030 67.595 ;
        RECT 109.170 67.515 119.300 67.625 ;
        RECT 109.170 67.495 114.715 67.515 ;
        RECT 109.170 67.455 114.215 67.495 ;
        RECT 109.170 67.180 109.340 67.455 ;
        RECT 108.725 67.010 109.340 67.180 ;
        RECT 109.825 66.885 119.300 67.055 ;
        RECT 109.825 66.170 109.995 66.885 ;
        RECT 111.290 66.255 119.300 66.425 ;
        RECT 109.105 65.170 110.105 66.170 ;
        RECT 111.290 65.660 111.460 66.255 ;
        RECT 110.830 65.490 111.460 65.660 ;
        RECT 111.010 65.450 111.460 65.490 ;
        RECT 112.000 65.625 119.300 65.795 ;
        RECT 112.000 64.755 112.170 65.625 ;
        RECT 109.980 64.585 112.170 64.755 ;
        RECT 112.610 64.995 119.300 65.165 ;
        RECT 102.270 64.325 102.800 64.440 ;
        RECT 93.520 63.425 94.750 63.595 ;
        RECT 95.070 63.980 100.645 64.150 ;
        RECT 101.080 64.025 102.800 64.325 ;
        RECT 109.980 64.225 110.150 64.585 ;
        RECT 93.520 62.930 93.690 63.425 ;
        RECT 92.725 61.930 93.725 62.930 ;
        RECT 95.070 62.655 95.240 63.980 ;
        RECT 95.895 63.350 100.645 63.520 ;
        RECT 96.295 62.930 96.465 63.350 ;
        RECT 101.080 63.270 101.410 64.025 ;
        RECT 102.270 63.910 102.800 64.025 ;
        RECT 109.105 63.640 110.150 64.225 ;
        RECT 112.610 63.905 112.780 64.995 ;
        RECT 111.215 63.835 112.780 63.905 ;
        RECT 111.035 63.735 112.780 63.835 ;
        RECT 113.230 64.365 119.300 64.535 ;
        RECT 111.035 63.665 111.565 63.735 ;
        RECT 109.105 63.225 110.105 63.640 ;
        RECT 113.230 63.350 113.400 64.365 ;
        RECT 112.170 63.180 113.400 63.350 ;
        RECT 113.720 63.735 119.300 63.905 ;
        RECT 94.645 62.620 95.240 62.655 ;
        RECT 94.465 62.485 95.240 62.620 ;
        RECT 94.465 62.450 94.995 62.485 ;
        RECT 95.880 61.930 96.880 62.930 ;
        RECT 112.170 62.685 112.340 63.180 ;
        RECT 111.375 61.685 112.375 62.685 ;
        RECT 113.720 62.410 113.890 63.735 ;
        RECT 114.550 63.105 119.300 63.275 ;
        RECT 114.945 62.685 115.115 63.105 ;
        RECT 119.735 63.025 120.065 69.180 ;
        RECT 113.295 62.375 113.890 62.410 ;
        RECT 113.115 62.240 113.890 62.375 ;
        RECT 113.115 62.205 113.645 62.240 ;
        RECT 114.530 61.685 115.530 62.685 ;
        RECT 105.380 56.575 106.045 56.745 ;
        RECT 69.880 54.530 70.180 54.795 ;
        RECT 69.880 54.230 70.425 54.530 ;
        RECT 72.505 54.470 73.035 55.000 ;
        RECT 56.440 53.300 56.970 53.830 ;
        RECT 50.020 53.150 50.190 53.155 ;
        RECT 50.020 52.980 55.800 53.150 ;
        RECT 70.125 52.985 70.425 54.230 ;
        RECT 82.260 53.155 82.560 55.215 ;
        RECT 104.480 55.170 105.480 55.640 ;
        RECT 105.875 55.630 106.045 56.575 ;
        RECT 106.730 56.050 107.730 57.050 ;
        RECT 108.385 56.575 109.165 56.745 ;
        RECT 107.465 55.840 107.635 56.050 ;
        RECT 107.465 55.670 108.670 55.840 ;
        RECT 105.875 55.460 107.135 55.630 ;
        RECT 106.965 55.205 107.135 55.460 ;
        RECT 104.480 55.000 106.620 55.170 ;
        RECT 106.965 55.035 108.175 55.205 ;
        RECT 104.480 54.640 105.480 55.000 ;
        RECT 106.450 54.645 106.620 55.000 ;
        RECT 106.450 54.475 107.650 54.645 ;
        RECT 107.480 54.025 107.650 54.475 ;
        RECT 108.005 54.535 108.175 55.035 ;
        RECT 108.500 55.050 108.670 55.670 ;
        RECT 108.995 55.570 109.165 56.575 ;
        RECT 109.730 56.635 110.730 57.050 ;
        RECT 109.730 56.050 110.800 56.635 ;
        RECT 108.995 55.400 110.330 55.570 ;
        RECT 108.500 54.880 109.850 55.050 ;
        RECT 108.005 54.365 109.390 54.535 ;
        RECT 82.260 52.985 82.590 53.155 ;
        RECT 50.020 52.540 50.190 52.980 ;
        RECT 49.560 51.540 50.560 52.540 ;
        RECT 70.010 52.455 70.540 52.985 ;
        RECT 82.165 52.455 82.695 52.985 ;
        RECT 104.145 52.965 105.145 53.965 ;
        RECT 107.480 53.855 108.875 54.025 ;
        RECT 105.935 53.500 107.000 53.670 ;
        RECT 106.830 53.430 107.000 53.500 ;
        RECT 106.830 53.260 108.375 53.430 ;
        RECT 104.815 52.620 104.985 52.965 ;
        RECT 49.275 50.470 50.365 50.800 ;
        RECT 58.190 50.755 59.080 51.645 ;
        RECT 62.320 51.090 63.050 51.095 ;
        RECT 62.140 51.080 63.050 51.090 ;
        RECT 62.140 50.925 69.740 51.080 ;
        RECT 62.140 50.920 62.670 50.925 ;
        RECT 62.950 50.910 69.740 50.925 ;
        RECT 49.275 46.260 49.605 50.470 ;
        RECT 49.835 50.430 50.365 50.470 ;
        RECT 50.030 49.790 50.200 50.430 ;
        RECT 59.575 50.170 60.575 50.650 ;
        RECT 59.575 50.000 69.740 50.170 ;
        RECT 50.030 49.620 55.800 49.790 ;
        RECT 59.575 49.650 60.575 50.000 ;
        RECT 62.320 49.270 63.180 49.275 ;
        RECT 62.140 49.260 63.180 49.270 ;
        RECT 62.140 49.105 69.740 49.260 ;
        RECT 62.140 49.100 62.670 49.105 ;
        RECT 62.950 49.090 69.740 49.105 ;
        RECT 59.575 48.350 60.575 48.765 ;
        RECT 56.460 47.730 56.990 48.260 ;
        RECT 59.575 48.180 69.740 48.350 ;
        RECT 59.575 47.765 60.575 48.180 ;
        RECT 62.320 47.450 63.160 47.455 ;
        RECT 62.140 47.440 63.160 47.450 ;
        RECT 62.140 47.285 69.740 47.440 ;
        RECT 62.140 47.280 62.670 47.285 ;
        RECT 62.950 47.270 69.740 47.285 ;
        RECT 59.575 46.530 60.575 46.940 ;
        RECT 50.020 46.510 50.190 46.530 ;
        RECT 50.020 46.340 55.800 46.510 ;
        RECT 59.575 46.360 69.740 46.530 ;
        RECT 50.020 45.915 50.190 46.340 ;
        RECT 59.575 45.940 60.575 46.360 ;
        RECT 35.430 43.995 36.680 45.245 ;
        RECT 49.560 44.915 50.560 45.915 ;
        RECT 62.150 45.615 62.680 45.630 ;
        RECT 62.950 45.615 69.740 45.620 ;
        RECT 62.150 45.460 69.740 45.615 ;
        RECT 62.330 45.450 69.740 45.460 ;
        RECT 62.330 45.445 63.050 45.450 ;
        RECT 59.575 44.710 60.575 45.065 ;
        RECT 59.575 44.540 69.740 44.710 ;
        RECT 42.000 44.130 42.530 44.300 ;
        RECT 35.805 43.670 36.105 43.995 ;
        RECT 35.805 40.060 36.135 43.670 ;
        RECT 42.175 43.590 42.345 44.130 ;
        RECT 46.575 44.125 47.105 44.295 ;
        RECT 36.610 43.420 42.380 43.590 ;
        RECT 42.175 43.410 42.345 43.420 ;
        RECT 45.930 42.270 46.260 43.670 ;
        RECT 46.750 43.590 46.920 44.125 ;
        RECT 59.575 44.065 60.575 44.540 ;
        RECT 62.150 43.795 62.680 43.810 ;
        RECT 62.950 43.795 69.740 43.800 ;
        RECT 62.150 43.640 69.740 43.795 ;
        RECT 62.330 43.630 69.740 43.640 ;
        RECT 62.330 43.625 63.100 43.630 ;
        RECT 46.735 43.420 52.505 43.590 ;
        RECT 46.750 43.405 46.920 43.420 ;
        RECT 45.175 42.155 46.260 42.270 ;
        RECT 59.575 42.890 60.575 43.245 ;
        RECT 59.575 42.720 69.740 42.890 ;
        RECT 59.575 42.245 60.575 42.720 ;
        RECT 43.160 41.570 43.690 42.100 ;
        RECT 45.075 41.985 46.260 42.155 ;
        RECT 62.330 41.985 63.195 41.995 ;
        RECT 45.175 41.940 46.260 41.985 ;
        RECT 36.610 40.140 42.380 40.310 ;
        RECT 37.945 39.685 38.115 40.140 ;
        RECT 45.930 40.060 46.260 41.940 ;
        RECT 62.150 41.980 63.195 41.985 ;
        RECT 62.150 41.825 69.740 41.980 ;
        RECT 62.150 41.815 62.680 41.825 ;
        RECT 62.950 41.810 69.740 41.825 ;
        RECT 53.220 41.155 53.750 41.685 ;
        RECT 59.575 41.070 60.575 41.505 ;
        RECT 59.575 40.900 69.740 41.070 ;
        RECT 59.575 40.505 60.575 40.900 ;
        RECT 46.735 40.140 52.505 40.310 ;
        RECT 62.140 40.160 63.185 40.175 ;
        RECT 46.755 39.695 46.925 40.140 ;
        RECT 62.140 40.005 69.740 40.160 ;
        RECT 62.950 39.990 69.740 40.005 ;
        RECT 37.485 38.685 38.485 39.685 ;
        RECT 46.295 38.695 47.295 39.695 ;
        RECT 59.575 39.250 60.575 39.670 ;
        RECT 59.575 39.080 69.740 39.250 ;
        RECT 59.575 38.670 60.575 39.080 ;
        RECT 35.430 37.265 36.680 38.515 ;
        RECT 62.415 38.355 62.610 38.470 ;
        RECT 62.415 38.350 63.145 38.355 ;
        RECT 62.150 38.340 63.145 38.350 ;
        RECT 62.150 38.185 69.740 38.340 ;
        RECT 62.150 38.180 62.680 38.185 ;
        RECT 62.950 38.170 69.740 38.185 ;
        RECT 70.155 38.090 70.485 52.455 ;
        RECT 72.830 50.620 73.440 51.290 ;
        RECT 73.830 50.615 74.360 50.795 ;
        RECT 82.260 50.700 82.590 52.455 ;
        RECT 104.815 52.450 107.780 52.620 ;
        RECT 105.075 51.495 106.930 51.500 ;
        RECT 104.895 51.330 106.930 51.495 ;
        RECT 104.895 51.325 105.425 51.330 ;
        RECT 75.070 50.615 81.860 50.620 ;
        RECT 73.830 50.450 81.860 50.615 ;
        RECT 82.260 50.490 82.605 50.700 ;
        RECT 73.830 50.445 75.250 50.450 ;
        RECT 73.830 50.265 74.360 50.445 ;
        RECT 71.110 49.335 72.110 49.765 ;
        RECT 75.070 49.335 81.860 49.340 ;
        RECT 71.110 49.170 81.860 49.335 ;
        RECT 71.110 49.165 75.245 49.170 ;
        RECT 71.110 48.765 72.110 49.165 ;
        RECT 73.755 48.055 74.285 48.230 ;
        RECT 75.070 48.055 81.860 48.060 ;
        RECT 73.755 47.890 81.860 48.055 ;
        RECT 73.755 47.885 75.140 47.890 ;
        RECT 73.755 47.700 74.285 47.885 ;
        RECT 71.050 46.775 72.050 47.195 ;
        RECT 75.070 46.775 81.860 46.780 ;
        RECT 71.050 46.610 81.860 46.775 ;
        RECT 71.050 46.605 75.140 46.610 ;
        RECT 71.050 46.195 72.050 46.605 ;
        RECT 73.750 45.495 74.280 45.675 ;
        RECT 75.070 45.495 81.860 45.500 ;
        RECT 73.750 45.330 81.860 45.495 ;
        RECT 73.750 45.325 75.140 45.330 ;
        RECT 73.750 45.145 74.280 45.325 ;
        RECT 71.160 44.215 72.160 44.690 ;
        RECT 75.070 44.215 81.860 44.220 ;
        RECT 71.160 44.050 81.860 44.215 ;
        RECT 71.160 44.045 75.140 44.050 ;
        RECT 71.160 43.690 72.160 44.045 ;
        RECT 73.790 42.935 74.320 43.110 ;
        RECT 75.070 42.935 81.860 42.940 ;
        RECT 73.790 42.770 81.860 42.935 ;
        RECT 73.790 42.765 75.140 42.770 ;
        RECT 73.790 42.580 74.320 42.765 ;
        RECT 71.160 41.655 72.160 42.080 ;
        RECT 75.070 41.655 81.860 41.660 ;
        RECT 71.160 41.490 81.860 41.655 ;
        RECT 71.160 41.485 75.140 41.490 ;
        RECT 71.160 41.080 72.160 41.485 ;
        RECT 73.765 40.375 74.295 40.550 ;
        RECT 75.070 40.375 81.860 40.380 ;
        RECT 73.765 40.210 81.860 40.375 ;
        RECT 73.765 40.205 75.140 40.210 ;
        RECT 73.765 40.020 74.295 40.205 ;
        RECT 71.160 39.095 72.160 39.595 ;
        RECT 75.070 39.095 81.860 39.100 ;
        RECT 71.160 38.930 81.860 39.095 ;
        RECT 71.160 38.925 75.140 38.930 ;
        RECT 71.160 38.595 72.160 38.925 ;
        RECT 42.020 37.470 42.550 37.640 ;
        RECT 46.575 37.495 47.105 37.665 ;
        RECT 75.070 37.650 81.860 37.820 ;
        RECT 35.810 36.975 36.130 37.265 ;
        RECT 35.805 33.365 36.135 36.975 ;
        RECT 42.195 36.895 42.365 37.470 ;
        RECT 36.610 36.725 42.380 36.895 ;
        RECT 43.130 34.865 43.660 35.395 ;
        RECT 45.930 35.225 46.260 36.975 ;
        RECT 46.750 36.895 46.920 37.495 ;
        RECT 74.240 36.945 74.770 37.125 ;
        RECT 75.830 36.945 76.000 37.650 ;
        RECT 82.275 37.570 82.605 50.490 ;
        RECT 106.760 50.545 106.930 51.330 ;
        RECT 107.610 51.175 107.780 52.450 ;
        RECT 108.205 51.805 108.375 53.260 ;
        RECT 108.705 52.435 108.875 53.855 ;
        RECT 109.220 53.065 109.390 54.365 ;
        RECT 109.680 53.695 109.850 54.880 ;
        RECT 110.160 54.325 110.330 55.400 ;
        RECT 110.630 54.955 110.800 56.050 ;
        RECT 112.270 55.585 112.970 56.745 ;
        RECT 111.715 55.415 118.505 55.585 ;
        RECT 110.630 54.785 118.505 54.955 ;
        RECT 110.160 54.155 118.505 54.325 ;
        RECT 109.680 53.525 118.505 53.695 ;
        RECT 109.220 52.895 118.505 53.065 ;
        RECT 108.705 52.265 118.505 52.435 ;
        RECT 108.205 51.635 118.505 51.805 ;
        RECT 107.610 51.005 118.505 51.175 ;
        RECT 118.920 50.550 119.250 55.665 ;
        RECT 106.760 50.375 118.505 50.545 ;
        RECT 104.145 49.915 105.145 50.345 ;
        RECT 104.145 49.745 118.505 49.915 ;
        RECT 118.920 49.850 120.625 50.550 ;
        RECT 104.145 49.345 105.145 49.745 ;
        RECT 106.600 49.115 118.505 49.285 ;
        RECT 106.600 48.220 106.770 49.115 ;
        RECT 105.075 48.215 106.770 48.220 ;
        RECT 104.895 48.050 106.770 48.215 ;
        RECT 107.490 48.655 111.880 48.665 ;
        RECT 107.490 48.495 118.505 48.655 ;
        RECT 104.895 48.045 105.425 48.050 ;
        RECT 107.490 47.355 107.660 48.495 ;
        RECT 111.715 48.485 118.505 48.495 ;
        RECT 106.695 47.185 107.660 47.355 ;
        RECT 108.100 47.855 118.505 48.025 ;
        RECT 106.695 47.100 106.865 47.185 ;
        RECT 104.560 46.930 106.865 47.100 ;
        RECT 104.560 46.595 104.730 46.930 ;
        RECT 108.100 46.680 108.270 47.855 ;
        RECT 104.145 45.595 105.145 46.595 ;
        RECT 107.305 46.510 108.270 46.680 ;
        RECT 108.625 47.225 118.505 47.395 ;
        RECT 107.305 46.175 107.475 46.510 ;
        RECT 105.935 46.005 107.475 46.175 ;
        RECT 108.625 46.060 108.795 47.225 ;
        RECT 107.845 45.890 108.795 46.060 ;
        RECT 109.210 46.595 118.505 46.765 ;
        RECT 107.845 45.060 108.015 45.890 ;
        RECT 109.210 45.480 109.380 46.595 ;
        RECT 104.820 44.505 105.820 44.990 ;
        RECT 106.855 44.890 108.015 45.060 ;
        RECT 108.385 45.310 109.380 45.480 ;
        RECT 109.700 45.965 118.505 46.135 ;
        RECT 106.855 44.505 107.025 44.890 ;
        RECT 104.820 44.335 107.025 44.505 ;
        RECT 108.385 44.480 108.555 45.310 ;
        RECT 109.700 44.870 109.870 45.965 ;
        RECT 104.820 43.990 105.820 44.335 ;
        RECT 107.520 44.310 108.555 44.480 ;
        RECT 108.905 44.700 109.870 44.870 ;
        RECT 110.260 45.335 118.505 45.505 ;
        RECT 107.520 44.045 107.690 44.310 ;
        RECT 106.430 43.875 107.690 44.045 ;
        RECT 108.905 43.995 109.075 44.700 ;
        RECT 110.260 44.230 110.430 45.335 ;
        RECT 106.430 43.045 106.600 43.875 ;
        RECT 108.070 43.825 109.075 43.995 ;
        RECT 109.415 44.060 110.430 44.230 ;
        RECT 110.920 44.705 118.505 44.875 ;
        RECT 108.070 43.500 108.240 43.825 ;
        RECT 105.935 42.875 106.600 43.045 ;
        RECT 106.115 42.865 106.600 42.875 ;
        RECT 107.230 42.915 108.240 43.500 ;
        RECT 109.415 43.045 109.585 44.060 ;
        RECT 110.920 43.540 111.090 44.705 ;
        RECT 111.715 44.075 118.505 44.245 ;
        RECT 112.525 44.070 112.705 44.075 ;
        RECT 109.015 43.020 109.585 43.045 ;
        RECT 107.230 42.500 108.230 42.915 ;
        RECT 108.835 42.875 109.585 43.020 ;
        RECT 109.960 42.970 111.090 43.540 ;
        RECT 112.535 43.275 112.705 44.070 ;
        RECT 118.920 43.995 119.250 49.850 ;
        RECT 112.355 43.105 112.885 43.275 ;
        RECT 108.835 42.850 109.365 42.875 ;
        RECT 109.960 42.540 110.960 42.970 ;
        RECT 110.945 40.510 111.475 41.040 ;
        RECT 46.735 36.725 52.505 36.895 ;
        RECT 74.240 36.775 76.000 36.945 ;
        RECT 74.240 36.595 74.770 36.775 ;
        RECT 56.035 35.350 56.565 35.680 ;
        RECT 45.175 35.190 46.260 35.225 ;
        RECT 45.075 35.020 46.260 35.190 ;
        RECT 45.175 34.895 46.260 35.020 ;
        RECT 36.610 33.445 42.380 33.615 ;
        RECT 37.595 32.980 37.765 33.445 ;
        RECT 45.930 33.365 46.260 34.895 ;
        RECT 53.240 34.820 53.770 35.350 ;
        RECT 56.235 33.995 56.565 35.350 ;
        RECT 57.135 34.460 58.135 35.460 ;
        RECT 71.030 34.875 71.920 35.765 ;
        RECT 56.835 33.995 57.165 34.040 ;
        RECT 56.235 33.665 57.165 33.995 ;
        RECT 57.635 33.960 57.805 34.460 ;
        RECT 57.580 33.790 64.370 33.960 ;
        RECT 46.735 33.445 52.505 33.615 ;
        RECT 46.740 32.990 46.910 33.445 ;
        RECT 35.430 31.170 36.680 32.420 ;
        RECT 37.135 31.980 38.135 32.980 ;
        RECT 46.280 31.990 47.280 32.990 ;
        RECT 56.835 32.800 57.165 33.665 ;
        RECT 64.740 33.100 65.350 33.770 ;
        RECT 70.285 33.745 70.615 34.215 ;
        RECT 71.465 34.135 71.635 34.875 ;
        RECT 71.030 33.965 77.820 34.135 ;
        RECT 69.215 33.685 70.615 33.745 ;
        RECT 69.115 33.515 70.615 33.685 ;
        RECT 69.215 33.415 70.615 33.515 ;
        RECT 57.580 32.880 64.370 33.050 ;
        RECT 70.285 32.975 70.615 33.415 ;
        RECT 71.030 33.055 77.820 33.225 ;
        RECT 78.790 33.220 79.400 33.890 ;
        RECT 57.595 32.415 57.765 32.880 ;
        RECT 41.980 31.355 42.510 31.525 ;
        RECT 35.815 30.860 36.135 31.170 ;
        RECT 35.805 27.250 36.135 30.860 ;
        RECT 42.155 30.780 42.325 31.355 ;
        RECT 47.765 31.335 48.295 31.505 ;
        RECT 57.135 31.415 58.135 32.415 ;
        RECT 71.675 32.335 71.845 33.055 ;
        RECT 71.495 31.805 72.025 32.335 ;
        RECT 36.610 30.610 42.380 30.780 ;
        RECT 43.130 28.775 43.660 29.305 ;
        RECT 45.930 28.985 46.260 30.860 ;
        RECT 47.940 30.780 48.110 31.335 ;
        RECT 46.735 30.610 52.505 30.780 ;
        RECT 45.075 28.655 46.260 28.985 ;
        RECT 53.240 28.795 53.770 29.325 ;
        RECT 36.610 27.330 42.380 27.500 ;
        RECT 37.595 26.865 37.765 27.330 ;
        RECT 45.930 27.250 46.260 28.655 ;
        RECT 46.775 27.500 46.945 27.510 ;
        RECT 46.735 27.330 52.505 27.500 ;
        RECT 46.775 26.895 46.945 27.330 ;
        RECT 35.600 24.800 36.850 26.050 ;
        RECT 37.135 25.865 38.135 26.865 ;
        RECT 46.315 25.895 47.315 26.895 ;
        RECT 61.695 26.415 61.865 27.085 ;
        RECT 42.020 24.930 42.550 25.100 ;
        RECT 47.765 24.930 48.295 25.100 ;
        RECT 35.820 24.455 36.120 24.800 ;
        RECT 35.805 20.845 36.135 24.455 ;
        RECT 42.195 24.375 42.365 24.930 ;
        RECT 36.610 24.205 42.380 24.375 ;
        RECT 45.930 22.900 46.260 24.455 ;
        RECT 47.940 24.375 48.110 24.930 ;
        RECT 46.735 24.205 52.505 24.375 ;
        RECT 61.695 23.995 61.865 25.875 ;
        RECT 86.760 25.205 86.930 27.085 ;
        RECT 45.175 22.830 46.260 22.900 ;
        RECT 43.130 22.300 43.660 22.830 ;
        RECT 45.075 22.660 46.260 22.830 ;
        RECT 45.175 22.570 46.260 22.660 ;
        RECT 36.610 21.085 42.380 21.095 ;
        RECT 36.605 20.925 42.380 21.085 ;
        RECT 36.605 20.470 36.775 20.925 ;
        RECT 45.930 20.845 46.260 22.570 ;
        RECT 53.240 22.450 53.770 22.980 ;
        RECT 61.695 21.575 61.865 23.455 ;
        RECT 86.760 22.785 86.930 24.665 ;
        RECT 86.760 21.575 86.930 22.245 ;
        RECT 46.730 21.095 46.900 21.105 ;
        RECT 46.730 20.925 52.505 21.095 ;
        RECT 46.730 20.490 46.900 20.925 ;
        RECT 36.145 19.470 37.145 20.470 ;
        RECT 46.270 19.490 47.270 20.490 ;
      LAYER met1 ;
        RECT 85.960 220.735 86.960 220.830 ;
        RECT 9.305 219.735 86.960 220.735 ;
        RECT 9.305 3.015 10.305 219.735 ;
        RECT 61.075 218.935 62.075 219.735 ;
        RECT 85.960 218.935 86.960 219.735 ;
        RECT 37.655 213.295 43.330 218.935 ;
        RECT 56.275 213.435 66.275 218.935 ;
        RECT 84.015 213.525 94.015 218.935 ;
        RECT 95.730 216.645 114.660 217.345 ;
        RECT 37.655 212.595 54.485 213.295 ;
        RECT 37.655 188.840 43.330 212.595 ;
        RECT 51.700 211.275 52.400 212.595 ;
        RECT 51.700 210.575 52.455 211.275 ;
        RECT 51.720 208.230 52.420 210.575 ;
        RECT 58.970 210.370 59.560 211.020 ;
        RECT 53.495 208.650 54.085 209.300 ;
        RECT 51.720 207.530 54.475 208.230 ;
        RECT 51.720 206.375 52.420 207.530 ;
        RECT 51.720 205.675 52.455 206.375 ;
        RECT 59.115 206.365 59.415 210.370 ;
        RECT 62.655 208.880 63.355 213.435 ;
        RECT 64.070 209.580 64.660 210.230 ;
        RECT 91.565 208.880 92.265 213.525 ;
        RECT 93.155 209.580 93.745 210.230 ;
        RECT 62.530 207.870 63.480 208.880 ;
        RECT 91.440 207.870 92.390 208.880 ;
        RECT 58.970 205.715 59.560 206.365 ;
        RECT 63.890 205.775 64.480 206.425 ;
        RECT 93.155 205.795 93.745 206.445 ;
        RECT 51.740 201.800 52.440 205.675 ;
        RECT 53.455 203.840 54.045 204.490 ;
        RECT 51.740 201.100 54.400 201.800 ;
        RECT 51.740 199.140 52.495 201.100 ;
        RECT 59.115 199.970 59.415 205.715 ;
        RECT 95.730 205.485 96.430 216.645 ;
        RECT 98.955 216.055 99.545 216.230 ;
        RECT 93.910 205.470 96.430 205.485 ;
        RECT 63.895 204.665 64.475 205.305 ;
        RECT 65.110 204.785 96.430 205.470 ;
        RECT 96.870 215.755 99.545 216.055 ;
        RECT 96.870 208.860 97.170 215.755 ;
        RECT 98.955 215.580 99.545 215.755 ;
        RECT 104.580 214.775 105.180 216.645 ;
        RECT 107.235 215.975 107.825 216.230 ;
        RECT 104.565 214.125 105.180 214.775 ;
        RECT 97.590 212.960 98.190 213.600 ;
        RECT 103.020 209.790 103.610 210.440 ;
        RECT 98.955 208.860 99.545 209.035 ;
        RECT 96.870 208.560 99.545 208.860 ;
        RECT 65.110 204.770 94.610 204.785 ;
        RECT 65.110 204.700 65.810 204.770 ;
        RECT 58.970 199.320 59.560 199.970 ;
        RECT 51.740 196.875 52.440 199.140 ;
        RECT 53.510 197.895 54.100 198.070 ;
        RECT 59.115 197.895 59.415 199.320 ;
        RECT 53.510 197.595 59.415 197.895 ;
        RECT 53.510 197.420 54.100 197.595 ;
        RECT 51.740 196.175 54.455 196.875 ;
        RECT 51.740 195.150 52.440 196.175 ;
        RECT 51.740 194.450 52.455 195.150 ;
        RECT 59.115 194.925 59.415 197.595 ;
        RECT 58.970 194.275 59.560 194.925 ;
        RECT 53.510 193.075 54.100 193.250 ;
        RECT 59.115 193.075 59.415 194.275 ;
        RECT 53.510 192.775 59.415 193.075 ;
        RECT 53.510 192.600 54.100 192.775 ;
        RECT 53.655 190.320 53.955 192.600 ;
        RECT 53.445 189.680 54.025 190.320 ;
        RECT 37.655 188.790 47.275 188.840 ;
        RECT 37.655 188.140 55.855 188.790 ;
        RECT 37.655 184.110 43.330 188.140 ;
        RECT 44.560 186.880 45.260 188.140 ;
        RECT 46.575 188.090 55.855 188.140 ;
        RECT 53.830 186.005 54.420 186.655 ;
        RECT 52.820 184.655 53.410 184.830 ;
        RECT 53.975 184.655 54.275 186.005 ;
        RECT 54.435 184.655 55.015 184.820 ;
        RECT 52.820 184.355 55.015 184.655 ;
        RECT 52.820 184.180 53.410 184.355 ;
        RECT 37.655 183.410 47.220 184.110 ;
        RECT 37.655 179.535 43.330 183.410 ;
        RECT 44.550 182.425 45.250 183.410 ;
        RECT 53.975 182.200 54.275 184.355 ;
        RECT 54.435 184.180 55.015 184.355 ;
        RECT 53.830 181.550 54.420 182.200 ;
        RECT 52.820 180.140 53.410 180.315 ;
        RECT 53.975 180.140 54.275 181.550 ;
        RECT 52.820 179.840 54.275 180.140 ;
        RECT 52.820 179.665 53.410 179.840 ;
        RECT 37.655 179.520 47.110 179.535 ;
        RECT 37.655 178.870 47.220 179.520 ;
        RECT 37.655 178.835 47.110 178.870 ;
        RECT 37.655 173.995 43.330 178.835 ;
        RECT 44.550 177.825 45.250 178.835 ;
        RECT 53.975 177.505 54.275 179.840 ;
        RECT 55.155 178.425 55.855 188.090 ;
        RECT 56.620 186.995 57.200 187.170 ;
        RECT 64.035 186.995 64.335 204.665 ;
        RECT 83.290 203.170 83.990 204.770 ;
        RECT 81.520 202.470 83.990 203.170 ;
        RECT 76.210 200.375 76.790 201.015 ;
        RECT 76.370 199.985 76.670 200.375 ;
        RECT 76.235 199.335 76.825 199.985 ;
        RECT 76.370 196.915 76.670 199.335 ;
        RECT 77.680 196.915 78.270 197.090 ;
        RECT 76.370 196.615 78.270 196.915 ;
        RECT 76.370 192.710 76.670 196.615 ;
        RECT 77.680 196.440 78.270 196.615 ;
        RECT 83.290 196.065 83.990 202.470 ;
        RECT 81.520 195.365 83.990 196.065 ;
        RECT 83.290 194.265 83.990 195.365 ;
        RECT 96.870 201.885 97.170 208.560 ;
        RECT 98.955 208.385 99.545 208.560 ;
        RECT 97.590 205.785 98.190 206.425 ;
        RECT 103.105 202.725 103.695 203.375 ;
        RECT 98.955 201.885 99.545 202.060 ;
        RECT 96.870 201.585 99.545 201.885 ;
        RECT 96.870 194.875 97.170 201.585 ;
        RECT 98.955 201.410 99.545 201.585 ;
        RECT 97.590 198.835 98.190 199.475 ;
        RECT 103.105 195.845 103.695 196.495 ;
        RECT 98.955 194.875 99.545 195.085 ;
        RECT 96.870 194.575 99.545 194.875 ;
        RECT 76.215 192.060 76.805 192.710 ;
        RECT 76.360 190.085 76.660 192.060 ;
        RECT 95.820 191.760 96.420 192.400 ;
        RECT 77.680 190.085 78.270 190.225 ;
        RECT 76.360 189.785 78.270 190.085 ;
        RECT 76.360 188.970 76.660 189.785 ;
        RECT 77.680 189.575 78.270 189.785 ;
        RECT 95.970 188.970 96.270 191.760 ;
        RECT 76.360 188.670 96.270 188.970 ;
        RECT 76.360 188.665 76.660 188.670 ;
        RECT 96.870 187.990 97.170 194.575 ;
        RECT 98.955 194.435 99.545 194.575 ;
        RECT 104.580 192.595 105.180 214.125 ;
        RECT 105.450 215.835 107.825 215.975 ;
        RECT 105.450 208.780 105.590 215.835 ;
        RECT 107.235 215.580 107.825 215.835 ;
        RECT 113.960 214.650 114.660 216.645 ;
        RECT 112.665 213.950 114.660 214.650 ;
        RECT 105.785 213.100 106.385 213.740 ;
        RECT 106.940 209.790 107.530 210.440 ;
        RECT 107.235 208.780 107.825 209.035 ;
        RECT 105.450 208.640 107.825 208.780 ;
        RECT 105.450 201.875 105.590 208.640 ;
        RECT 107.235 208.385 107.825 208.640 ;
        RECT 113.960 207.885 114.660 213.950 ;
        RECT 112.665 207.185 114.660 207.885 ;
        RECT 105.785 206.020 106.385 206.660 ;
        RECT 107.025 202.725 107.615 203.375 ;
        RECT 107.235 201.875 107.825 202.130 ;
        RECT 105.450 201.735 107.825 201.875 ;
        RECT 105.450 194.895 105.590 201.735 ;
        RECT 107.235 201.480 107.825 201.735 ;
        RECT 112.610 200.690 113.310 200.750 ;
        RECT 113.960 200.690 114.660 207.185 ;
        RECT 112.610 199.990 114.660 200.690 ;
        RECT 105.785 199.150 106.385 199.790 ;
        RECT 107.025 195.845 107.615 196.495 ;
        RECT 107.235 194.895 107.825 195.150 ;
        RECT 105.450 194.755 107.825 194.895 ;
        RECT 97.590 191.810 98.190 192.450 ;
        RECT 103.105 188.685 103.695 189.335 ;
        RECT 105.450 187.990 105.590 194.755 ;
        RECT 107.235 194.500 107.825 194.755 ;
        RECT 113.960 193.270 114.660 199.990 ;
        RECT 120.150 193.270 124.655 218.935 ;
        RECT 112.665 192.570 124.655 193.270 ;
        RECT 105.785 191.810 106.385 192.450 ;
        RECT 107.025 188.685 107.615 189.335 ;
        RECT 96.870 187.690 119.730 187.990 ;
        RECT 56.620 186.695 64.335 186.995 ;
        RECT 56.620 186.530 57.200 186.695 ;
        RECT 58.515 184.060 58.745 185.920 ;
        RECT 118.850 185.720 119.080 185.920 ;
        RECT 119.430 185.720 119.730 187.690 ;
        RECT 118.850 185.580 119.730 185.720 ;
        RECT 118.850 185.270 119.080 185.580 ;
        RECT 58.515 181.640 58.745 183.500 ;
        RECT 118.850 182.850 119.080 184.710 ;
        RECT 58.515 179.220 58.745 181.080 ;
        RECT 118.850 180.430 119.080 182.290 ;
        RECT 120.150 179.870 124.655 192.570 ;
        RECT 118.850 179.220 124.655 179.870 ;
        RECT 55.155 177.725 88.690 178.425 ;
        RECT 53.830 176.855 54.420 177.505 ;
        RECT 52.820 175.535 53.410 175.715 ;
        RECT 53.975 175.535 54.275 176.855 ;
        RECT 52.820 175.235 54.275 175.535 ;
        RECT 52.820 175.065 53.410 175.235 ;
        RECT 37.655 173.950 46.710 173.995 ;
        RECT 37.655 173.300 47.135 173.950 ;
        RECT 37.655 173.295 46.710 173.300 ;
        RECT 37.655 169.515 43.330 173.295 ;
        RECT 44.550 172.280 45.250 173.295 ;
        RECT 53.975 171.795 54.275 175.235 ;
        RECT 87.990 174.570 88.690 177.725 ;
        RECT 104.880 176.225 113.735 176.925 ;
        RECT 89.220 175.565 89.810 176.215 ;
        RECT 87.865 173.560 88.815 174.570 ;
        RECT 104.880 174.300 105.580 176.225 ;
        RECT 107.055 176.055 107.645 176.225 ;
        RECT 91.160 173.600 105.580 174.300 ;
        RECT 113.035 174.965 113.735 176.225 ;
        RECT 120.150 174.965 124.655 179.220 ;
        RECT 113.035 174.265 124.655 174.965 ;
        RECT 53.805 171.145 54.395 171.795 ;
        RECT 37.655 168.815 47.190 169.515 ;
        RECT 52.585 169.465 53.175 170.115 ;
        RECT 37.655 164.860 43.330 168.815 ;
        RECT 44.630 167.665 45.330 168.815 ;
        RECT 53.975 167.485 54.275 171.145 ;
        RECT 53.835 166.835 54.425 167.485 ;
        RECT 46.490 164.860 47.190 164.925 ;
        RECT 37.655 164.160 47.190 164.860 ;
        RECT 52.520 164.830 53.110 165.480 ;
        RECT 21.385 148.680 23.625 148.745 ;
        RECT 37.655 148.680 43.330 164.160 ;
        RECT 44.550 163.175 45.250 164.160 ;
        RECT 53.975 162.885 54.275 166.835 ;
        RECT 87.990 164.610 88.690 173.560 ;
        RECT 89.245 171.595 89.835 172.245 ;
        RECT 89.235 165.505 89.825 166.155 ;
        RECT 87.955 163.600 88.905 164.610 ;
        RECT 92.270 164.380 92.970 173.600 ;
        RECT 105.755 172.745 106.355 173.385 ;
        RECT 107.275 170.790 107.865 170.880 ;
        RECT 105.155 170.490 107.865 170.790 ;
        RECT 93.960 165.970 94.550 166.185 ;
        RECT 105.155 165.970 105.455 170.490 ;
        RECT 107.275 170.230 107.865 170.490 ;
        RECT 107.000 169.480 107.700 169.535 ;
        RECT 107.000 168.780 113.725 169.480 ;
        RECT 113.025 168.410 113.725 168.780 ;
        RECT 120.150 168.410 124.655 174.265 ;
        RECT 113.025 167.735 124.655 168.410 ;
        RECT 113.080 167.710 124.655 167.735 ;
        RECT 93.960 165.670 105.455 165.970 ;
        RECT 105.755 165.955 106.355 166.595 ;
        RECT 93.960 165.535 94.550 165.670 ;
        RECT 91.170 163.680 92.970 164.380 ;
        RECT 105.155 163.575 105.455 165.670 ;
        RECT 107.275 163.575 107.865 163.750 ;
        RECT 105.155 163.275 107.865 163.575 ;
        RECT 107.275 163.100 107.865 163.275 ;
        RECT 53.815 162.235 54.405 162.885 ;
        RECT 86.105 162.095 86.720 162.100 ;
        RECT 86.070 160.730 86.720 162.095 ;
        RECT 89.245 161.605 89.835 162.255 ;
        RECT 52.525 160.080 53.115 160.730 ;
        RECT 55.465 160.030 113.610 160.730 ;
        RECT 86.070 160.020 86.720 160.030 ;
        RECT 112.910 158.260 113.610 160.030 ;
        RECT 45.875 156.400 46.105 158.260 ;
        RECT 110.880 157.610 113.610 158.260 ;
        RECT 45.875 153.980 46.105 155.840 ;
        RECT 110.880 155.190 111.110 157.050 ;
        RECT 45.875 151.560 46.105 153.420 ;
        RECT 110.880 152.770 111.110 154.630 ;
        RECT 45.875 149.140 46.105 151.000 ;
        RECT 110.880 150.350 111.110 152.210 ;
        RECT 21.385 146.680 43.330 148.680 ;
        RECT 45.875 146.720 46.105 148.580 ;
        RECT 110.880 147.930 111.110 149.790 ;
        RECT 21.385 146.545 23.625 146.680 ;
        RECT 37.655 138.900 43.330 146.680 ;
        RECT 45.875 144.300 46.105 146.160 ;
        RECT 110.880 145.510 111.110 147.370 ;
        RECT 112.910 145.835 113.610 157.610 ;
        RECT 120.150 147.680 124.655 167.710 ;
        RECT 138.235 147.680 140.475 147.760 ;
        RECT 45.875 141.880 46.105 143.740 ;
        RECT 110.880 143.090 111.110 144.950 ;
        RECT 45.875 139.460 46.105 141.320 ;
        RECT 110.880 140.670 111.110 142.530 ;
        RECT 110.880 139.460 112.180 140.110 ;
        RECT 111.530 138.900 112.180 139.460 ;
        RECT 37.655 138.250 112.180 138.900 ;
        RECT 37.655 137.935 43.330 138.250 ;
        RECT 112.655 137.935 117.655 145.835 ;
        RECT 120.150 145.680 140.475 147.680 ;
        RECT 120.150 137.935 124.655 145.680 ;
        RECT 138.235 145.560 140.475 145.680 ;
        RECT 114.645 115.410 115.645 137.935 ;
        RECT 14.115 114.410 115.645 115.410 ;
        RECT 14.115 4.490 15.115 114.410 ;
        RECT 28.775 88.185 34.885 110.400 ;
        RECT 44.040 108.150 44.940 108.310 ;
        RECT 53.025 108.160 53.925 108.320 ;
        RECT 63.260 108.160 64.160 108.320 ;
        RECT 44.020 107.510 44.960 108.150 ;
        RECT 53.005 107.520 53.945 108.160 ;
        RECT 63.240 107.520 64.180 108.160 ;
        RECT 71.665 108.135 72.245 108.775 ;
        RECT 76.765 108.685 77.665 108.845 ;
        RECT 44.040 107.350 44.940 107.510 ;
        RECT 53.025 107.360 53.925 107.520 ;
        RECT 63.260 107.360 64.160 107.520 ;
        RECT 42.285 105.635 43.185 105.795 ;
        RECT 42.265 104.995 43.205 105.635 ;
        RECT 59.500 105.490 60.400 105.650 ;
        RECT 69.525 105.490 70.425 105.650 ;
        RECT 42.285 104.835 43.185 104.995 ;
        RECT 49.735 104.700 50.325 105.350 ;
        RECT 59.480 104.850 60.420 105.490 ;
        RECT 69.505 104.850 70.445 105.490 ;
        RECT 71.775 105.145 71.915 108.135 ;
        RECT 76.745 108.045 77.685 108.685 ;
        RECT 76.765 107.885 77.665 108.045 ;
        RECT 79.950 106.570 80.530 106.755 ;
        RECT 124.150 106.570 129.030 110.400 ;
        RECT 79.905 105.870 129.030 106.570 ;
        RECT 43.965 101.165 44.965 102.165 ;
        RECT 44.040 99.300 44.940 99.460 ;
        RECT 44.020 98.660 44.960 99.300 ;
        RECT 44.040 98.500 44.940 98.660 ;
        RECT 49.975 96.475 50.115 104.700 ;
        RECT 59.500 104.690 60.400 104.850 ;
        RECT 69.525 104.690 70.425 104.850 ;
        RECT 71.535 104.495 72.125 105.145 ;
        RECT 80.355 104.865 80.935 105.060 ;
        RECT 80.355 104.725 81.305 104.865 ;
        RECT 52.175 102.735 52.765 103.385 ;
        RECT 49.960 96.275 50.115 96.475 ;
        RECT 42.285 95.840 43.185 96.000 ;
        RECT 42.265 95.200 43.205 95.840 ;
        RECT 49.960 95.240 50.100 96.275 ;
        RECT 42.285 95.040 43.185 95.200 ;
        RECT 49.755 94.590 50.345 95.240 ;
        RECT 43.965 91.255 44.965 92.255 ;
        RECT 35.365 88.185 35.945 88.435 ;
        RECT 28.775 88.045 35.945 88.185 ;
        RECT 44.040 88.080 44.940 88.240 ;
        RECT 28.775 57.190 34.885 88.045 ;
        RECT 35.365 87.795 35.945 88.045 ;
        RECT 44.020 87.440 44.960 88.080 ;
        RECT 44.040 87.280 44.940 87.440 ;
        RECT 42.285 86.480 43.185 86.640 ;
        RECT 42.265 85.840 43.205 86.480 ;
        RECT 42.285 85.680 43.185 85.840 ;
        RECT 49.960 85.165 50.100 94.590 ;
        RECT 52.400 93.455 52.540 102.735 ;
        RECT 62.335 102.705 62.925 103.355 ;
        RECT 52.950 101.200 53.950 102.200 ;
        RECT 62.555 99.025 62.695 102.705 ;
        RECT 63.445 101.140 64.445 102.140 ;
        RECT 71.775 101.810 71.915 104.495 ;
        RECT 80.355 104.420 80.935 104.725 ;
        RECT 81.165 103.920 81.305 104.725 ;
        RECT 81.110 103.270 81.340 103.920 ;
        RECT 72.385 101.810 73.335 102.180 ;
        RECT 71.775 101.670 73.335 101.810 ;
        RECT 77.415 101.775 78.315 101.935 ;
        RECT 71.775 99.025 71.915 101.670 ;
        RECT 72.385 101.170 73.335 101.670 ;
        RECT 77.395 101.135 78.335 101.775 ;
        RECT 77.415 100.975 78.315 101.135 ;
        RECT 81.110 100.850 81.340 102.710 ;
        RECT 121.945 102.060 122.175 103.920 ;
        RECT 62.555 98.885 71.915 99.025 ;
        RECT 53.025 98.200 53.925 98.360 ;
        RECT 53.005 97.560 53.945 98.200 ;
        RECT 53.025 97.400 53.925 97.560 ;
        RECT 62.555 97.160 62.695 98.885 ;
        RECT 63.260 98.220 64.160 98.380 ;
        RECT 63.240 97.580 64.180 98.220 ;
        RECT 63.260 97.420 64.160 97.580 ;
        RECT 62.335 96.510 62.925 97.160 ;
        RECT 59.500 95.140 60.400 95.300 ;
        RECT 59.480 94.500 60.420 95.140 ;
        RECT 59.500 94.340 60.400 94.500 ;
        RECT 52.175 92.805 52.765 93.455 ;
        RECT 49.735 84.515 50.325 85.165 ;
        RECT 43.965 81.100 44.965 82.100 ;
        RECT 44.040 79.005 44.940 79.165 ;
        RECT 44.020 78.365 44.960 79.005 ;
        RECT 44.040 78.205 44.940 78.365 ;
        RECT 41.680 75.995 42.580 76.155 ;
        RECT 41.660 75.355 42.600 75.995 ;
        RECT 49.960 75.965 50.100 84.515 ;
        RECT 52.400 83.405 52.540 92.805 ;
        RECT 52.950 91.290 53.950 92.290 ;
        RECT 53.025 88.430 53.925 88.590 ;
        RECT 53.005 87.790 53.945 88.430 ;
        RECT 53.025 87.630 53.925 87.790 ;
        RECT 62.555 87.155 62.695 96.510 ;
        RECT 69.525 95.140 70.425 95.300 ;
        RECT 71.775 95.180 71.915 98.885 ;
        RECT 76.690 98.685 77.590 98.845 ;
        RECT 76.670 98.045 77.610 98.685 ;
        RECT 81.110 98.430 81.340 100.290 ;
        RECT 121.945 99.640 122.175 101.500 ;
        RECT 124.150 99.085 129.030 105.870 ;
        RECT 122.070 99.080 129.030 99.085 ;
        RECT 121.945 98.430 129.030 99.080 ;
        RECT 122.070 98.385 129.030 98.430 ;
        RECT 76.690 97.885 77.590 98.045 ;
        RECT 124.150 97.885 129.030 98.385 ;
        RECT 120.190 97.185 129.030 97.885 ;
        RECT 91.515 96.710 110.825 96.850 ;
        RECT 69.505 94.500 70.445 95.140 ;
        RECT 71.555 94.530 72.145 95.180 ;
        RECT 91.515 95.120 91.655 96.710 ;
        RECT 110.685 95.715 110.825 96.710 ;
        RECT 91.400 94.850 91.990 95.120 ;
        RECT 84.235 94.710 91.990 94.850 ;
        RECT 69.525 94.340 70.425 94.500 ;
        RECT 63.445 91.245 64.445 92.245 ;
        RECT 71.775 91.800 71.915 94.530 ;
        RECT 72.385 91.800 73.335 92.280 ;
        RECT 77.415 92.255 78.315 92.415 ;
        RECT 71.775 91.660 73.335 91.800 ;
        RECT 63.260 88.555 64.160 88.715 ;
        RECT 63.240 87.915 64.180 88.555 ;
        RECT 63.260 87.755 64.160 87.915 ;
        RECT 62.335 86.505 62.925 87.155 ;
        RECT 59.500 85.120 60.400 85.280 ;
        RECT 59.480 84.480 60.420 85.120 ;
        RECT 59.500 84.320 60.400 84.480 ;
        RECT 52.175 82.755 52.765 83.405 ;
        RECT 52.390 79.815 52.530 82.755 ;
        RECT 52.950 81.275 53.950 82.275 ;
        RECT 62.560 79.815 62.700 86.505 ;
        RECT 69.525 85.280 70.425 85.440 ;
        RECT 71.775 85.420 71.915 91.660 ;
        RECT 72.385 91.270 73.335 91.660 ;
        RECT 77.395 91.615 78.335 92.255 ;
        RECT 77.415 91.455 78.315 91.615 ;
        RECT 76.690 88.855 77.590 89.015 ;
        RECT 76.670 88.215 77.610 88.855 ;
        RECT 76.690 88.055 77.590 88.215 ;
        RECT 69.505 84.640 70.445 85.280 ;
        RECT 71.495 84.770 72.085 85.420 ;
        RECT 69.525 84.480 70.425 84.640 ;
        RECT 71.775 83.515 71.915 84.770 ;
        RECT 71.760 83.375 71.915 83.515 ;
        RECT 63.445 81.390 64.445 82.390 ;
        RECT 52.390 79.675 62.700 79.815 ;
        RECT 52.390 77.985 52.530 79.675 ;
        RECT 53.025 78.995 53.925 79.155 ;
        RECT 53.005 78.355 53.945 78.995 ;
        RECT 53.025 78.195 53.925 78.355 ;
        RECT 52.175 77.335 52.765 77.985 ;
        RECT 62.560 77.890 62.700 79.675 ;
        RECT 63.260 79.040 64.160 79.200 ;
        RECT 63.240 78.400 64.180 79.040 ;
        RECT 63.260 78.240 64.160 78.400 ;
        RECT 62.335 77.240 62.925 77.890 ;
        RECT 59.500 76.185 60.400 76.345 ;
        RECT 49.755 75.700 50.345 75.965 ;
        RECT 50.530 75.700 51.110 75.950 ;
        RECT 49.755 75.560 51.110 75.700 ;
        RECT 41.680 75.195 42.580 75.355 ;
        RECT 49.755 75.315 50.345 75.560 ;
        RECT 50.530 75.310 51.110 75.560 ;
        RECT 59.480 75.545 60.420 76.185 ;
        RECT 69.525 75.955 70.425 76.115 ;
        RECT 59.500 75.385 60.400 75.545 ;
        RECT 69.505 75.315 70.445 75.955 ;
        RECT 71.775 75.720 71.915 83.375 ;
        RECT 72.490 81.540 73.490 82.540 ;
        RECT 77.380 81.900 78.280 82.060 ;
        RECT 77.360 81.260 78.300 81.900 ;
        RECT 77.380 81.100 78.280 81.260 ;
        RECT 76.850 78.730 77.750 78.890 ;
        RECT 76.830 78.090 77.770 78.730 ;
        RECT 76.850 77.930 77.750 78.090 ;
        RECT 84.235 76.105 84.375 94.710 ;
        RECT 91.400 94.470 91.990 94.710 ;
        RECT 94.635 94.465 95.635 95.465 ;
        RECT 96.140 95.090 97.040 95.250 ;
        RECT 96.120 94.450 97.060 95.090 ;
        RECT 110.435 95.065 111.025 95.715 ;
        RECT 112.965 94.465 113.965 95.465 ;
        RECT 114.470 95.090 115.370 95.250 ;
        RECT 114.450 94.450 115.390 95.090 ;
        RECT 96.140 94.290 97.040 94.450 ;
        RECT 114.470 94.290 115.370 94.450 ;
        RECT 94.210 93.840 95.110 94.000 ;
        RECT 112.540 93.840 113.440 94.000 ;
        RECT 92.730 92.740 93.730 93.740 ;
        RECT 94.190 93.200 95.130 93.840 ;
        RECT 94.210 93.040 95.110 93.200 ;
        RECT 91.700 91.175 92.700 92.175 ;
        RECT 93.160 92.170 94.060 92.330 ;
        RECT 93.140 91.530 94.080 92.170 ;
        RECT 102.765 92.055 103.765 93.055 ;
        RECT 111.060 92.740 112.060 93.740 ;
        RECT 112.520 93.200 113.460 93.840 ;
        RECT 112.540 93.040 113.440 93.200 ;
        RECT 93.160 91.370 94.060 91.530 ;
        RECT 110.030 91.175 111.030 92.175 ;
        RECT 111.490 92.170 112.390 92.330 ;
        RECT 111.470 91.530 112.410 92.170 ;
        RECT 111.490 91.370 112.390 91.530 ;
        RECT 87.845 89.775 88.745 89.935 ;
        RECT 87.825 89.135 88.765 89.775 ;
        RECT 89.350 89.670 90.350 90.670 ;
        RECT 91.045 90.590 91.945 90.750 ;
        RECT 91.025 89.950 91.965 90.590 ;
        RECT 91.045 89.790 91.945 89.950 ;
        RECT 106.175 89.775 107.075 89.935 ;
        RECT 106.155 89.135 107.095 89.775 ;
        RECT 107.680 89.670 108.680 90.670 ;
        RECT 109.375 90.590 110.275 90.750 ;
        RECT 109.355 89.950 110.295 90.590 ;
        RECT 109.375 89.790 110.275 89.950 ;
        RECT 87.845 88.975 88.745 89.135 ;
        RECT 106.175 88.975 107.075 89.135 ;
        RECT 86.135 87.510 87.135 88.510 ;
        RECT 87.845 87.415 88.745 87.575 ;
        RECT 104.465 87.530 105.465 88.530 ;
        RECT 124.150 88.485 129.030 97.185 ;
        RECT 120.055 87.785 129.030 88.485 ;
        RECT 106.175 87.415 107.075 87.575 ;
        RECT 87.825 86.775 88.765 87.415 ;
        RECT 106.155 86.775 107.095 87.415 ;
        RECT 87.845 86.615 88.745 86.775 ;
        RECT 106.175 86.615 107.075 86.775 ;
        RECT 88.670 85.130 89.670 86.130 ;
        RECT 90.180 85.950 91.080 86.110 ;
        RECT 90.160 85.310 91.100 85.950 ;
        RECT 90.180 85.150 91.080 85.310 ;
        RECT 107.000 85.130 108.000 86.130 ;
        RECT 108.510 85.950 109.410 86.110 ;
        RECT 108.490 85.310 109.430 85.950 ;
        RECT 108.510 85.150 109.410 85.310 ;
        RECT 90.745 83.705 91.745 84.705 ;
        RECT 92.285 84.430 93.185 84.590 ;
        RECT 92.265 83.790 93.205 84.430 ;
        RECT 92.285 83.630 93.185 83.790 ;
        RECT 109.075 83.705 110.075 84.705 ;
        RECT 110.615 84.430 111.515 84.590 ;
        RECT 110.595 83.790 111.535 84.430 ;
        RECT 110.615 83.630 111.515 83.790 ;
        RECT 90.745 81.760 91.745 82.760 ;
        RECT 92.490 82.605 93.390 82.765 ;
        RECT 92.470 81.965 93.410 82.605 ;
        RECT 92.490 81.805 93.390 81.965 ;
        RECT 109.075 81.760 110.075 82.760 ;
        RECT 110.820 82.605 111.720 82.765 ;
        RECT 110.800 81.965 111.740 82.605 ;
        RECT 110.820 81.805 111.720 81.965 ;
        RECT 93.015 80.220 94.015 81.220 ;
        RECT 94.570 81.145 95.470 81.305 ;
        RECT 94.550 80.505 95.490 81.145 ;
        RECT 94.570 80.345 95.470 80.505 ;
        RECT 96.170 80.220 97.170 81.220 ;
        RECT 111.345 80.220 112.345 81.220 ;
        RECT 112.900 81.145 113.800 81.305 ;
        RECT 112.880 80.505 113.820 81.145 ;
        RECT 112.900 80.345 113.800 80.505 ;
        RECT 114.500 80.220 115.500 81.220 ;
        RECT 91.265 77.870 110.105 78.010 ;
        RECT 91.265 76.735 91.405 77.870 ;
        RECT 91.090 76.105 91.680 76.735 ;
        RECT 94.395 76.175 95.395 77.175 ;
        RECT 95.850 76.800 96.750 76.960 ;
        RECT 95.830 76.160 96.770 76.800 ;
        RECT 109.965 76.360 110.105 77.870 ;
        RECT 84.235 76.085 91.680 76.105 ;
        RECT 84.235 75.965 91.405 76.085 ;
        RECT 95.850 76.000 96.750 76.160 ;
        RECT 69.525 75.155 70.425 75.315 ;
        RECT 71.515 75.070 72.105 75.720 ;
        RECT 43.965 72.095 44.965 73.095 ;
        RECT 52.950 72.070 53.950 73.070 ;
        RECT 63.445 72.215 64.445 73.215 ;
        RECT 72.085 71.915 73.085 72.915 ;
        RECT 77.510 72.380 78.410 72.540 ;
        RECT 77.490 71.740 78.430 72.380 ;
        RECT 77.510 71.580 78.410 71.740 ;
        RECT 49.725 71.000 50.625 71.160 ;
        RECT 49.705 70.360 50.645 71.000 ;
        RECT 49.725 70.200 50.625 70.360 ;
        RECT 56.450 68.415 57.030 69.055 ;
        RECT 56.635 67.710 56.775 68.415 ;
        RECT 72.540 68.245 73.120 68.495 ;
        RECT 73.800 68.245 74.390 68.500 ;
        RECT 61.720 68.030 62.620 68.190 ;
        RECT 72.540 68.105 74.390 68.245 ;
        RECT 56.410 67.060 57.000 67.710 ;
        RECT 61.700 67.390 62.640 68.030 ;
        RECT 72.540 67.855 73.120 68.105 ;
        RECT 73.800 67.850 74.390 68.105 ;
        RECT 61.720 67.230 62.620 67.390 ;
        RECT 49.560 64.895 50.560 65.895 ;
        RECT 49.725 64.460 50.625 64.620 ;
        RECT 49.705 63.820 50.645 64.460 ;
        RECT 49.725 63.660 50.625 63.820 ;
        RECT 56.650 62.375 56.790 67.060 ;
        RECT 61.720 66.210 62.620 66.370 ;
        RECT 61.700 65.570 62.640 66.210 ;
        RECT 74.025 65.985 74.165 67.850 ;
        RECT 61.720 65.410 62.620 65.570 ;
        RECT 73.800 65.335 74.390 65.985 ;
        RECT 61.720 64.390 62.620 64.550 ;
        RECT 61.700 63.750 62.640 64.390 ;
        RECT 61.720 63.590 62.620 63.750 ;
        RECT 74.025 63.380 74.165 65.335 ;
        RECT 61.730 62.575 62.630 62.735 ;
        RECT 73.800 62.730 74.390 63.380 ;
        RECT 56.430 61.725 57.020 62.375 ;
        RECT 61.710 61.935 62.650 62.575 ;
        RECT 61.730 61.775 62.630 61.935 ;
        RECT 46.010 58.790 46.590 59.020 ;
        RECT 43.320 58.650 46.590 58.790 ;
        RECT 28.775 57.175 35.880 57.190 ;
        RECT 28.775 56.535 36.170 57.175 ;
        RECT 28.775 56.490 35.880 56.535 ;
        RECT 28.775 46.515 34.885 56.490 ;
        RECT 28.775 45.815 36.170 46.515 ;
        RECT 28.775 44.960 34.885 45.815 ;
        RECT 35.400 44.960 36.710 45.305 ;
        RECT 28.775 44.260 36.710 44.960 ;
        RECT 41.815 44.535 42.715 44.695 ;
        RECT 28.775 38.380 34.885 44.260 ;
        RECT 35.400 43.935 36.710 44.260 ;
        RECT 41.795 43.895 42.735 44.535 ;
        RECT 41.815 43.735 42.715 43.895 ;
        RECT 43.320 42.160 43.460 58.650 ;
        RECT 46.010 58.380 46.590 58.650 ;
        RECT 49.560 58.205 50.560 59.205 ;
        RECT 49.725 57.765 50.625 57.925 ;
        RECT 49.705 57.125 50.645 57.765 ;
        RECT 49.725 56.965 50.625 57.125 ;
        RECT 56.635 53.890 56.775 61.725 ;
        RECT 61.730 60.750 62.630 60.910 ;
        RECT 74.025 60.850 74.165 62.730 ;
        RECT 61.710 60.110 62.650 60.750 ;
        RECT 73.800 60.200 74.390 60.850 ;
        RECT 61.730 59.950 62.630 60.110 ;
        RECT 61.730 58.925 62.630 59.085 ;
        RECT 61.710 58.285 62.650 58.925 ;
        RECT 61.730 58.125 62.630 58.285 ;
        RECT 74.025 58.205 74.165 60.200 ;
        RECT 73.800 57.555 74.390 58.205 ;
        RECT 61.720 57.115 62.620 57.275 ;
        RECT 61.700 56.475 62.640 57.115 ;
        RECT 61.720 56.315 62.620 56.475 ;
        RECT 74.025 55.730 74.165 57.555 ;
        RECT 59.425 55.290 60.325 55.450 ;
        RECT 61.730 55.290 62.630 55.450 ;
        RECT 59.405 54.650 60.345 55.290 ;
        RECT 61.710 54.650 62.650 55.290 ;
        RECT 73.800 55.080 74.390 55.730 ;
        RECT 71.220 54.805 71.800 55.070 ;
        RECT 72.475 54.805 73.065 55.060 ;
        RECT 71.220 54.665 73.065 54.805 ;
        RECT 59.425 54.490 60.325 54.650 ;
        RECT 61.730 54.490 62.630 54.650 ;
        RECT 71.220 54.430 71.800 54.665 ;
        RECT 72.475 54.410 73.065 54.665 ;
        RECT 84.235 54.335 84.375 75.965 ;
        RECT 109.740 75.710 110.330 76.360 ;
        RECT 112.995 75.930 113.995 76.930 ;
        RECT 114.500 76.555 115.400 76.715 ;
        RECT 114.480 75.915 115.420 76.555 ;
        RECT 114.500 75.755 115.400 75.915 ;
        RECT 93.920 75.550 94.820 75.710 ;
        RECT 92.440 74.450 93.440 75.450 ;
        RECT 93.900 74.910 94.840 75.550 ;
        RECT 112.570 75.305 113.470 75.465 ;
        RECT 93.920 74.750 94.820 74.910 ;
        RECT 111.090 74.205 112.090 75.205 ;
        RECT 112.550 74.665 113.490 75.305 ;
        RECT 112.570 74.505 113.470 74.665 ;
        RECT 91.410 72.885 92.410 73.885 ;
        RECT 92.870 73.880 93.770 74.040 ;
        RECT 92.850 73.240 93.790 73.880 ;
        RECT 92.870 73.080 93.770 73.240 ;
        RECT 110.060 72.640 111.060 73.640 ;
        RECT 111.520 73.635 112.420 73.795 ;
        RECT 111.500 72.995 112.440 73.635 ;
        RECT 111.520 72.835 112.420 72.995 ;
        RECT 87.555 71.485 88.455 71.645 ;
        RECT 87.535 70.845 88.475 71.485 ;
        RECT 89.060 71.380 90.060 72.380 ;
        RECT 90.755 72.300 91.655 72.460 ;
        RECT 90.735 71.660 91.675 72.300 ;
        RECT 90.755 71.500 91.655 71.660 ;
        RECT 106.205 71.240 107.105 71.400 ;
        RECT 87.555 70.685 88.455 70.845 ;
        RECT 106.185 70.600 107.125 71.240 ;
        RECT 107.710 71.135 108.710 72.135 ;
        RECT 109.405 72.055 110.305 72.215 ;
        RECT 109.385 71.415 110.325 72.055 ;
        RECT 109.405 71.255 110.305 71.415 ;
        RECT 106.205 70.440 107.105 70.600 ;
        RECT 85.845 69.240 86.845 70.240 ;
        RECT 87.555 69.125 88.455 69.285 ;
        RECT 87.535 68.485 88.475 69.125 ;
        RECT 104.495 69.010 105.495 70.010 ;
        RECT 124.150 69.880 129.030 87.785 ;
        RECT 120.340 69.180 129.030 69.880 ;
        RECT 106.205 68.880 107.105 69.040 ;
        RECT 87.555 68.325 88.455 68.485 ;
        RECT 106.185 68.240 107.125 68.880 ;
        RECT 106.205 68.080 107.105 68.240 ;
        RECT 88.380 66.840 89.380 67.840 ;
        RECT 89.890 67.660 90.790 67.820 ;
        RECT 89.870 67.020 90.810 67.660 ;
        RECT 89.890 66.860 90.790 67.020 ;
        RECT 107.030 66.595 108.030 67.595 ;
        RECT 108.540 67.415 109.440 67.575 ;
        RECT 108.520 66.775 109.460 67.415 ;
        RECT 108.540 66.615 109.440 66.775 ;
        RECT 90.455 65.415 91.455 66.415 ;
        RECT 91.995 66.140 92.895 66.300 ;
        RECT 91.975 65.500 92.915 66.140 ;
        RECT 91.995 65.340 92.895 65.500 ;
        RECT 109.105 65.170 110.105 66.170 ;
        RECT 110.645 65.895 111.545 66.055 ;
        RECT 110.625 65.255 111.565 65.895 ;
        RECT 110.645 65.095 111.545 65.255 ;
        RECT 90.455 63.470 91.455 64.470 ;
        RECT 92.200 64.315 93.100 64.475 ;
        RECT 92.180 63.675 93.120 64.315 ;
        RECT 102.240 64.125 102.830 64.500 ;
        RECT 92.200 63.515 93.100 63.675 ;
        RECT 92.725 61.930 93.725 62.930 ;
        RECT 94.280 62.855 95.180 63.015 ;
        RECT 94.260 62.215 95.200 62.855 ;
        RECT 94.280 62.055 95.180 62.215 ;
        RECT 95.880 61.930 96.880 62.930 ;
        RECT 102.185 60.035 102.885 64.125 ;
        RECT 109.105 63.225 110.105 64.225 ;
        RECT 110.850 64.070 111.750 64.230 ;
        RECT 110.830 63.430 111.770 64.070 ;
        RECT 110.850 63.270 111.750 63.430 ;
        RECT 111.375 61.685 112.375 62.685 ;
        RECT 112.930 62.610 113.830 62.770 ;
        RECT 112.910 61.970 113.850 62.610 ;
        RECT 112.930 61.810 113.830 61.970 ;
        RECT 114.530 61.685 115.530 62.685 ;
        RECT 124.150 60.035 129.030 69.180 ;
        RECT 102.185 59.335 129.030 60.035 ;
        RECT 102.215 58.665 102.915 59.335 ;
        RECT 73.935 54.195 84.375 54.335 ;
        RECT 99.730 57.965 102.915 58.665 ;
        RECT 56.410 53.240 57.000 53.890 ;
        RECT 73.935 53.855 74.075 54.195 ;
        RECT 58.510 53.715 74.075 53.855 ;
        RECT 49.560 51.540 50.560 52.540 ;
        RECT 49.650 50.835 50.550 50.995 ;
        RECT 49.630 50.195 50.570 50.835 ;
        RECT 49.650 50.035 50.550 50.195 ;
        RECT 56.650 48.320 56.790 53.240 ;
        RECT 58.510 51.705 58.650 53.715 ;
        RECT 99.730 53.070 100.430 57.965 ;
        RECT 105.195 56.980 106.095 57.140 ;
        RECT 105.175 56.340 106.115 56.980 ;
        RECT 105.195 56.180 106.095 56.340 ;
        RECT 106.730 56.050 107.730 57.050 ;
        RECT 108.200 56.980 109.100 57.140 ;
        RECT 108.180 56.340 109.120 56.980 ;
        RECT 108.200 56.180 109.100 56.340 ;
        RECT 109.730 56.050 110.730 57.050 ;
        RECT 112.170 56.980 113.070 57.140 ;
        RECT 112.150 56.340 113.090 56.980 ;
        RECT 112.170 56.180 113.070 56.340 ;
        RECT 104.480 54.640 105.480 55.640 ;
        RECT 69.980 52.370 100.430 53.070 ;
        RECT 104.145 52.965 105.145 53.965 ;
        RECT 105.750 53.905 106.650 54.065 ;
        RECT 105.730 53.265 106.670 53.905 ;
        RECT 105.750 53.105 106.650 53.265 ;
        RECT 58.160 50.695 59.110 51.705 ;
        RECT 61.955 51.325 62.855 51.485 ;
        RECT 58.565 49.145 58.705 50.695 ;
        RECT 61.935 50.685 62.875 51.325 ;
        RECT 71.220 51.025 71.800 51.320 ;
        RECT 72.840 51.025 73.430 51.280 ;
        RECT 71.220 50.885 73.430 51.025 ;
        RECT 59.575 49.650 60.575 50.650 ;
        RECT 61.955 50.525 62.855 50.685 ;
        RECT 71.220 50.680 71.800 50.885 ;
        RECT 72.840 50.630 73.430 50.885 ;
        RECT 73.745 50.880 74.445 52.370 ;
        RECT 104.710 51.730 105.610 51.890 ;
        RECT 104.690 51.090 105.630 51.730 ;
        RECT 104.710 50.930 105.610 51.090 ;
        RECT 73.685 50.600 74.445 50.880 ;
        RECT 73.685 50.460 74.560 50.600 ;
        RECT 124.150 50.590 129.030 59.335 ;
        RECT 73.685 50.180 74.445 50.460 ;
        RECT 61.955 49.505 62.855 49.665 ;
        RECT 58.270 48.505 58.850 49.145 ;
        RECT 61.935 48.865 62.875 49.505 ;
        RECT 56.430 47.670 57.020 48.320 ;
        RECT 59.575 47.765 60.575 48.765 ;
        RECT 61.955 48.705 62.855 48.865 ;
        RECT 71.110 48.765 72.110 49.765 ;
        RECT 73.950 48.290 74.090 50.180 ;
        RECT 104.145 49.345 105.145 50.345 ;
        RECT 119.980 49.890 129.030 50.590 ;
        RECT 104.710 48.450 105.610 48.610 ;
        RECT 61.955 47.685 62.855 47.845 ;
        RECT 61.935 47.045 62.875 47.685 ;
        RECT 73.725 47.640 74.315 48.290 ;
        RECT 104.690 47.810 105.630 48.450 ;
        RECT 104.710 47.650 105.610 47.810 ;
        RECT 59.575 45.940 60.575 46.940 ;
        RECT 61.955 46.885 62.855 47.045 ;
        RECT 71.050 46.195 72.050 47.195 ;
        RECT 49.560 44.915 50.560 45.915 ;
        RECT 61.965 45.865 62.865 46.025 ;
        RECT 61.945 45.225 62.885 45.865 ;
        RECT 73.945 45.735 74.085 47.640 ;
        RECT 61.965 45.065 62.865 45.225 ;
        RECT 73.720 45.085 74.310 45.735 ;
        RECT 104.145 45.595 105.145 46.595 ;
        RECT 105.750 46.410 106.650 46.570 ;
        RECT 105.730 45.770 106.670 46.410 ;
        RECT 105.750 45.610 106.650 45.770 ;
        RECT 46.390 44.530 47.290 44.690 ;
        RECT 46.370 43.890 47.310 44.530 ;
        RECT 59.575 44.065 60.575 45.065 ;
        RECT 61.965 44.045 62.865 44.205 ;
        RECT 46.390 43.730 47.290 43.890 ;
        RECT 61.945 43.405 62.885 44.045 ;
        RECT 71.160 43.690 72.160 44.690 ;
        RECT 61.965 43.245 62.865 43.405 ;
        RECT 44.890 42.390 45.790 42.550 ;
        RECT 43.130 41.510 43.720 42.160 ;
        RECT 44.870 41.750 45.810 42.390 ;
        RECT 59.575 42.245 60.575 43.245 ;
        RECT 73.985 43.170 74.125 45.085 ;
        RECT 104.820 43.990 105.820 44.990 ;
        RECT 105.750 43.280 106.650 43.440 ;
        RECT 73.760 42.520 74.350 43.170 ;
        RECT 105.730 42.640 106.670 43.280 ;
        RECT 61.965 42.220 62.865 42.380 ;
        RECT 44.890 41.590 45.790 41.750 ;
        RECT 37.485 38.685 38.485 39.685 ;
        RECT 35.400 38.380 36.710 38.575 ;
        RECT 28.775 37.680 36.710 38.380 ;
        RECT 41.835 37.875 42.735 38.035 ;
        RECT 28.775 31.885 34.885 37.680 ;
        RECT 35.400 37.205 36.710 37.680 ;
        RECT 41.815 37.235 42.755 37.875 ;
        RECT 41.835 37.075 42.735 37.235 ;
        RECT 43.320 36.085 43.460 41.510 ;
        RECT 53.190 41.095 53.780 41.745 ;
        RECT 61.945 41.580 62.885 42.220 ;
        RECT 46.295 38.695 47.295 39.695 ;
        RECT 46.390 37.900 47.290 38.060 ;
        RECT 46.370 37.260 47.310 37.900 ;
        RECT 46.390 37.100 47.290 37.260 ;
        RECT 53.430 36.085 53.570 41.095 ;
        RECT 59.575 40.505 60.575 41.505 ;
        RECT 61.965 41.420 62.865 41.580 ;
        RECT 71.160 41.080 72.160 42.080 ;
        RECT 73.960 40.610 74.100 42.520 ;
        RECT 105.750 42.480 106.650 42.640 ;
        RECT 107.230 42.500 108.230 43.500 ;
        RECT 108.650 43.255 109.550 43.415 ;
        RECT 108.630 42.615 109.570 43.255 ;
        RECT 108.650 42.455 109.550 42.615 ;
        RECT 109.960 42.540 110.960 43.540 ;
        RECT 112.170 43.510 113.070 43.670 ;
        RECT 112.150 42.870 113.090 43.510 ;
        RECT 124.150 43.490 129.030 49.890 ;
        RECT 123.875 43.440 129.030 43.490 ;
        RECT 112.170 42.710 113.070 42.870 ;
        RECT 123.510 42.800 129.030 43.440 ;
        RECT 123.875 42.790 129.030 42.800 ;
        RECT 61.955 40.410 62.855 40.570 ;
        RECT 61.935 39.770 62.875 40.410 ;
        RECT 73.735 39.960 74.325 40.610 ;
        RECT 110.915 40.450 111.505 41.100 ;
        RECT 59.575 38.670 60.575 39.670 ;
        RECT 61.955 39.610 62.855 39.770 ;
        RECT 61.965 38.585 62.865 38.745 ;
        RECT 71.160 38.595 72.160 39.595 ;
        RECT 61.945 37.945 62.885 38.585 ;
        RECT 61.965 37.785 62.865 37.945 ;
        RECT 71.255 37.560 71.835 37.730 ;
        RECT 68.225 37.260 72.850 37.560 ;
        RECT 43.320 35.940 43.465 36.085 ;
        RECT 53.430 35.940 53.575 36.085 ;
        RECT 43.325 35.455 43.465 35.940 ;
        RECT 43.100 34.805 43.690 35.455 ;
        RECT 44.890 35.425 45.790 35.585 ;
        RECT 35.400 31.885 36.710 32.480 ;
        RECT 37.135 31.980 38.135 32.980 ;
        RECT 28.775 31.185 36.710 31.885 ;
        RECT 41.795 31.760 42.695 31.920 ;
        RECT 21.385 29.655 23.625 29.665 ;
        RECT 28.775 29.655 34.885 31.185 ;
        RECT 35.400 31.110 36.710 31.185 ;
        RECT 41.775 31.120 42.715 31.760 ;
        RECT 41.795 30.960 42.695 31.120 ;
        RECT 21.385 27.655 34.885 29.655 ;
        RECT 43.325 29.365 43.465 34.805 ;
        RECT 44.870 34.785 45.810 35.425 ;
        RECT 53.435 35.410 53.575 35.940 ;
        RECT 55.850 35.835 56.750 35.995 ;
        RECT 44.890 34.625 45.790 34.785 ;
        RECT 53.210 34.760 53.800 35.410 ;
        RECT 55.830 35.195 56.770 35.835 ;
        RECT 55.850 35.035 56.750 35.195 ;
        RECT 46.280 31.990 47.280 32.990 ;
        RECT 47.580 31.740 48.480 31.900 ;
        RECT 47.560 31.100 48.500 31.740 ;
        RECT 47.580 30.940 48.480 31.100 ;
        RECT 53.435 29.385 53.575 34.760 ;
        RECT 57.135 34.460 58.135 35.460 ;
        RECT 64.750 33.700 65.340 33.760 ;
        RECT 64.750 33.110 65.480 33.700 ;
        RECT 57.135 31.415 58.135 32.415 ;
        RECT 43.100 28.715 43.690 29.365 ;
        RECT 44.890 29.140 45.790 29.300 ;
        RECT 21.385 27.465 23.625 27.655 ;
        RECT 28.775 25.660 34.885 27.655 ;
        RECT 35.570 25.660 36.880 26.110 ;
        RECT 37.135 25.865 38.135 26.865 ;
        RECT 28.775 24.960 36.880 25.660 ;
        RECT 41.835 25.335 42.735 25.495 ;
        RECT 28.775 17.075 34.885 24.960 ;
        RECT 35.570 24.740 36.880 24.960 ;
        RECT 41.815 24.695 42.755 25.335 ;
        RECT 41.835 24.535 42.735 24.695 ;
        RECT 43.325 22.890 43.465 28.715 ;
        RECT 44.870 28.500 45.810 29.140 ;
        RECT 53.210 28.735 53.800 29.385 ;
        RECT 44.890 28.340 45.790 28.500 ;
        RECT 46.315 25.895 47.315 26.895 ;
        RECT 47.580 25.335 48.480 25.495 ;
        RECT 47.560 24.695 48.500 25.335 ;
        RECT 47.580 24.535 48.480 24.695 ;
        RECT 44.890 23.065 45.790 23.225 ;
        RECT 43.100 22.240 43.690 22.890 ;
        RECT 44.870 22.425 45.810 23.065 ;
        RECT 53.435 23.040 53.575 28.735 ;
        RECT 55.060 26.425 61.895 27.075 ;
        RECT 44.890 22.265 45.790 22.425 ;
        RECT 53.210 22.390 53.800 23.040 ;
        RECT 36.145 19.470 37.145 20.470 ;
        RECT 43.325 18.005 43.465 22.240 ;
        RECT 46.270 19.490 47.270 20.490 ;
        RECT 53.435 18.005 53.575 22.390 ;
        RECT 43.325 17.865 53.575 18.005 ;
        RECT 55.060 17.075 55.710 26.425 ;
        RECT 61.665 24.005 61.895 25.865 ;
        RECT 61.665 21.585 61.895 23.445 ;
        RECT 28.775 16.425 55.710 17.075 ;
        RECT 28.775 10.610 34.885 16.425 ;
        RECT 64.780 15.875 65.480 33.110 ;
        RECT 68.225 32.210 68.525 37.260 ;
        RECT 71.255 37.090 71.835 37.260 ;
        RECT 72.550 36.350 72.850 37.260 ;
        RECT 73.905 36.930 74.045 39.960 ;
        RECT 111.140 39.620 111.280 40.450 ;
        RECT 110.840 38.980 111.420 39.620 ;
        RECT 74.210 36.930 74.800 37.185 ;
        RECT 73.905 36.790 74.800 36.930 ;
        RECT 74.210 36.535 74.800 36.790 ;
        RECT 71.000 34.815 71.950 35.825 ;
        RECT 72.485 35.710 73.065 36.350 ;
        RECT 68.930 33.920 69.830 34.080 ;
        RECT 68.910 33.280 69.850 33.920 ;
        RECT 68.930 33.120 69.830 33.280 ;
        RECT 71.465 32.210 72.055 32.395 ;
        RECT 68.225 31.910 72.055 32.210 ;
        RECT 71.465 31.745 72.055 31.910 ;
        RECT 55.505 10.595 65.505 15.875 ;
        RECT 78.735 15.690 79.435 33.950 ;
        RECT 86.730 25.215 86.960 27.075 ;
        RECT 86.730 22.795 86.960 24.655 ;
        RECT 86.730 21.585 87.940 22.235 ;
        RECT 87.290 18.445 87.940 21.585 ;
        RECT 95.355 18.445 96.355 18.620 ;
        RECT 87.290 17.795 96.355 18.445 ;
        RECT 87.290 15.860 87.940 17.795 ;
        RECT 95.355 17.620 96.355 17.795 ;
        RECT 124.150 16.850 129.030 42.790 ;
        RECT 138.235 16.850 140.475 16.930 ;
        RECT 69.445 10.615 79.445 15.690 ;
        RECT 86.410 10.620 96.410 15.860 ;
        RECT 124.150 14.850 140.475 16.850 ;
        RECT 63.860 6.225 64.860 10.595 ;
        RECT 77.650 8.130 78.650 10.615 ;
        RECT 91.800 10.070 92.800 10.620 ;
        RECT 124.150 10.610 129.030 14.850 ;
        RECT 138.235 14.730 140.475 14.850 ;
        RECT 138.715 10.070 139.995 10.210 ;
        RECT 91.800 9.070 139.995 10.070 ;
        RECT 138.715 8.970 139.995 9.070 ;
        RECT 77.650 8.000 129.095 8.130 ;
        RECT 77.650 7.130 129.665 8.000 ;
        RECT 128.385 6.760 129.665 7.130 ;
        RECT 63.860 6.080 106.850 6.225 ;
        RECT 63.860 5.225 107.730 6.080 ;
        RECT 106.450 4.840 107.730 5.225 ;
        RECT 14.115 4.415 85.085 4.490 ;
        RECT 14.115 3.865 85.390 4.415 ;
        RECT 14.155 3.490 85.390 3.865 ;
        RECT 84.110 3.175 85.390 3.490 ;
        RECT 9.305 2.875 62.350 3.015 ;
        RECT 9.305 2.015 63.215 2.875 ;
        RECT 61.935 1.635 63.215 2.015 ;
      LAYER met2 ;
        RECT 97.525 212.895 98.255 213.665 ;
        RECT 105.720 213.035 106.450 213.805 ;
        RECT 103.025 210.335 103.605 210.435 ;
        RECT 106.945 210.335 107.525 210.435 ;
        RECT 64.075 210.055 64.655 210.225 ;
        RECT 93.160 210.055 93.740 210.225 ;
        RECT 103.025 210.195 107.525 210.335 ;
        RECT 64.075 209.755 95.270 210.055 ;
        RECT 103.025 209.795 103.605 210.195 ;
        RECT 64.075 209.585 64.655 209.755 ;
        RECT 93.160 209.585 93.740 209.755 ;
        RECT 53.500 209.095 54.080 209.295 ;
        RECT 53.500 208.795 60.805 209.095 ;
        RECT 53.500 208.655 54.080 208.795 ;
        RECT 53.460 204.255 54.040 204.485 ;
        RECT 60.505 204.255 60.805 208.795 ;
        RECT 63.895 206.270 64.475 206.420 ;
        RECT 93.160 206.270 93.740 206.440 ;
        RECT 63.895 205.970 93.740 206.270 ;
        RECT 63.895 205.780 64.475 205.970 ;
        RECT 93.160 205.800 93.740 205.970 ;
        RECT 64.035 205.305 64.335 205.780 ;
        RECT 63.895 204.665 64.475 205.305 ;
        RECT 53.460 203.955 76.610 204.255 ;
        RECT 53.460 203.845 54.040 203.955 ;
        RECT 76.310 201.015 76.610 203.955 ;
        RECT 76.210 200.375 76.790 201.015 ;
        RECT 53.170 189.415 54.300 190.585 ;
        RECT 56.620 186.530 57.200 187.170 ;
        RECT 54.435 184.650 55.015 184.820 ;
        RECT 56.765 184.650 57.065 186.530 ;
        RECT 54.435 184.350 57.065 184.650 ;
        RECT 54.435 184.180 55.015 184.350 ;
        RECT 89.225 176.040 89.805 176.210 ;
        RECT 89.225 176.000 93.525 176.040 ;
        RECT 94.970 176.000 95.270 209.755 ;
        RECT 97.525 205.720 98.255 206.490 ;
        RECT 103.110 203.120 103.690 203.370 ;
        RECT 105.255 203.120 105.395 210.195 ;
        RECT 106.945 209.795 107.525 210.195 ;
        RECT 105.720 205.955 106.450 206.725 ;
        RECT 107.030 203.120 107.610 203.370 ;
        RECT 103.110 202.980 107.610 203.120 ;
        RECT 103.110 202.730 103.690 202.980 ;
        RECT 97.525 198.770 98.255 199.540 ;
        RECT 103.110 196.240 103.690 196.490 ;
        RECT 105.255 196.240 105.395 202.980 ;
        RECT 107.030 202.730 107.610 202.980 ;
        RECT 105.720 199.085 106.450 199.855 ;
        RECT 107.030 196.240 107.610 196.490 ;
        RECT 103.110 196.100 107.610 196.240 ;
        RECT 103.110 195.850 103.690 196.100 ;
        RECT 95.755 191.695 96.485 192.465 ;
        RECT 97.525 191.745 98.255 192.515 ;
        RECT 97.525 189.080 98.255 189.485 ;
        RECT 103.110 189.080 103.690 189.330 ;
        RECT 105.255 189.080 105.395 196.100 ;
        RECT 107.030 195.850 107.610 196.100 ;
        RECT 105.720 191.745 106.450 192.515 ;
        RECT 107.030 189.080 107.610 189.330 ;
        RECT 97.525 188.940 107.610 189.080 ;
        RECT 97.525 188.715 98.255 188.940 ;
        RECT 103.110 188.690 103.690 188.940 ;
        RECT 107.030 188.690 107.610 188.940 ;
        RECT 89.225 175.740 95.270 176.000 ;
        RECT 89.225 175.570 89.805 175.740 ;
        RECT 93.225 175.700 95.270 175.740 ;
        RECT 89.250 172.025 89.830 172.240 ;
        RECT 86.210 171.725 89.830 172.025 ;
        RECT 52.735 170.150 53.435 170.155 ;
        RECT 52.505 169.450 55.225 170.150 ;
        RECT 52.525 165.470 53.105 165.475 ;
        RECT 54.525 165.470 55.225 169.450 ;
        RECT 52.525 164.835 55.225 165.470 ;
        RECT 52.565 164.770 55.225 164.835 ;
        RECT 52.530 160.710 53.425 160.725 ;
        RECT 54.525 160.710 55.225 164.770 ;
        RECT 86.210 162.095 86.510 171.725 ;
        RECT 89.250 171.600 89.830 171.725 ;
        RECT 89.240 165.980 89.820 166.150 ;
        RECT 93.225 165.980 93.525 175.700 ;
        RECT 105.690 172.680 106.420 173.450 ;
        RECT 93.965 165.980 94.545 166.180 ;
        RECT 89.240 165.680 94.545 165.980 ;
        RECT 105.690 165.890 106.420 166.660 ;
        RECT 89.240 165.510 89.820 165.680 ;
        RECT 93.965 165.540 94.545 165.680 ;
        RECT 86.105 162.080 86.685 162.095 ;
        RECT 89.250 162.080 89.830 162.250 ;
        RECT 86.105 161.780 89.830 162.080 ;
        RECT 86.105 161.455 86.685 161.780 ;
        RECT 89.250 161.610 89.830 161.780 ;
        RECT 55.405 160.710 56.105 160.725 ;
        RECT 52.470 160.010 56.105 160.710 ;
        RECT 21.320 146.480 23.690 148.810 ;
        RECT 138.170 145.495 140.540 147.825 ;
        RECT 52.145 109.035 81.005 109.175 ;
        RECT 44.040 108.120 44.940 108.310 ;
        RECT 41.585 107.420 44.940 108.120 ;
        RECT 41.585 105.795 42.285 107.420 ;
        RECT 44.040 107.350 44.940 107.420 ;
        RECT 52.145 107.910 52.285 109.035 ;
        RECT 53.025 107.910 53.925 108.320 ;
        RECT 52.145 107.770 53.925 107.910 ;
        RECT 41.585 104.835 43.185 105.795 ;
        RECT 41.585 99.445 42.285 104.835 ;
        RECT 43.900 101.080 45.030 102.250 ;
        RECT 44.040 99.445 44.940 99.460 ;
        RECT 41.585 98.745 44.940 99.445 ;
        RECT 41.585 96.000 42.285 98.745 ;
        RECT 43.910 98.710 44.940 98.745 ;
        RECT 44.040 98.500 44.940 98.710 ;
        RECT 52.145 97.860 52.285 107.770 ;
        RECT 53.025 107.360 53.925 107.770 ;
        RECT 62.330 107.910 62.470 109.035 ;
        RECT 63.260 107.910 64.160 108.320 ;
        RECT 71.590 108.070 72.320 108.840 ;
        RECT 76.765 108.785 77.665 108.845 ;
        RECT 76.765 108.085 79.720 108.785 ;
        RECT 62.330 107.770 64.160 107.910 ;
        RECT 76.765 107.885 77.665 108.085 ;
        RECT 59.500 105.520 60.400 105.650 ;
        RECT 59.480 104.690 60.400 105.520 ;
        RECT 52.885 101.115 54.015 102.285 ;
        RECT 53.025 97.860 53.925 98.360 ;
        RECT 52.135 97.720 53.925 97.860 ;
        RECT 41.585 95.040 43.185 96.000 ;
        RECT 35.365 88.425 35.945 88.435 ;
        RECT 41.585 88.425 42.285 95.040 ;
        RECT 43.900 91.170 45.030 92.340 ;
        RECT 35.365 88.240 44.490 88.425 ;
        RECT 35.365 87.795 44.940 88.240 ;
        RECT 52.145 88.180 52.285 97.720 ;
        RECT 53.025 97.400 53.925 97.720 ;
        RECT 59.480 95.300 60.180 104.690 ;
        RECT 62.330 97.880 62.470 107.770 ;
        RECT 63.260 107.360 64.160 107.770 ;
        RECT 79.020 106.830 79.720 108.085 ;
        RECT 79.020 106.130 80.590 106.830 ;
        RECT 69.525 104.690 70.425 105.650 ;
        RECT 63.380 101.055 64.510 102.225 ;
        RECT 63.260 97.880 64.160 98.380 ;
        RECT 62.330 97.740 64.160 97.880 ;
        RECT 59.480 94.340 60.400 95.300 ;
        RECT 52.885 91.205 54.015 92.375 ;
        RECT 53.025 88.180 53.925 88.590 ;
        RECT 52.135 88.040 53.925 88.180 ;
        RECT 35.655 87.725 44.940 87.795 ;
        RECT 41.585 86.640 42.285 87.725 ;
        RECT 44.040 87.280 44.940 87.725 ;
        RECT 41.585 85.680 43.185 86.640 ;
        RECT 41.585 78.995 42.285 85.680 ;
        RECT 43.900 81.015 45.030 82.185 ;
        RECT 44.040 78.995 44.940 79.165 ;
        RECT 41.585 78.295 44.940 78.995 ;
        RECT 52.145 78.715 52.285 88.040 ;
        RECT 53.025 87.630 53.925 88.040 ;
        RECT 59.480 85.280 60.180 94.340 ;
        RECT 62.330 88.305 62.470 97.740 ;
        RECT 63.260 97.420 64.160 97.740 ;
        RECT 69.625 95.300 70.325 104.690 ;
        RECT 77.415 101.805 78.315 101.935 ;
        RECT 77.400 100.975 78.315 101.805 ;
        RECT 77.400 100.835 78.100 100.975 ;
        RECT 79.020 100.835 79.720 106.130 ;
        RECT 79.890 106.115 80.590 106.130 ;
        RECT 80.865 105.060 81.005 109.035 ;
        RECT 80.355 104.670 81.005 105.060 ;
        RECT 80.355 104.420 80.935 104.670 ;
        RECT 76.760 100.135 79.720 100.835 ;
        RECT 76.760 98.845 77.460 100.135 ;
        RECT 76.690 97.885 77.590 98.845 ;
        RECT 69.525 94.340 70.425 95.300 ;
        RECT 63.380 91.160 64.510 92.330 ;
        RECT 63.260 88.305 64.160 88.715 ;
        RECT 62.330 88.165 64.160 88.305 ;
        RECT 59.480 84.320 60.400 85.280 ;
        RECT 52.885 81.190 54.015 82.360 ;
        RECT 53.025 78.715 53.925 79.155 ;
        RECT 52.145 78.575 53.925 78.715 ;
        RECT 41.585 76.155 42.285 78.295 ;
        RECT 44.040 78.205 44.940 78.295 ;
        RECT 53.025 78.195 53.925 78.575 ;
        RECT 59.480 76.345 60.180 84.320 ;
        RECT 62.330 78.745 62.470 88.165 ;
        RECT 63.260 87.755 64.160 88.165 ;
        RECT 69.625 85.440 70.325 94.340 ;
        RECT 77.415 91.455 78.315 92.415 ;
        RECT 77.515 90.560 78.215 91.455 ;
        RECT 79.020 90.560 79.720 100.135 ;
        RECT 120.125 97.150 120.855 97.920 ;
        RECT 94.115 96.010 114.970 96.150 ;
        RECT 94.115 94.000 94.255 96.010 ;
        RECT 94.570 94.380 95.700 95.550 ;
        RECT 96.460 95.250 96.600 96.010 ;
        RECT 96.140 94.290 97.040 95.250 ;
        RECT 92.665 92.655 93.795 93.825 ;
        RECT 94.115 93.450 95.110 94.000 ;
        RECT 94.210 93.040 95.110 93.450 ;
        RECT 76.735 89.860 79.720 90.560 ;
        RECT 88.225 91.435 91.140 91.575 ;
        RECT 88.225 89.935 88.365 91.435 ;
        RECT 76.735 89.015 77.435 89.860 ;
        RECT 76.690 88.055 77.590 89.015 ;
        RECT 69.525 84.480 70.425 85.440 ;
        RECT 63.380 81.305 64.510 82.475 ;
        RECT 63.260 78.745 64.160 79.200 ;
        RECT 62.330 78.605 64.160 78.745 ;
        RECT 63.260 78.240 64.160 78.605 ;
        RECT 41.585 75.325 42.580 76.155 ;
        RECT 41.680 75.195 42.580 75.325 ;
        RECT 50.455 75.245 51.185 76.015 ;
        RECT 59.480 75.385 60.400 76.345 ;
        RECT 69.625 76.115 70.325 84.480 ;
        RECT 72.425 81.455 73.555 82.625 ;
        RECT 77.380 81.100 78.280 82.060 ;
        RECT 77.555 80.365 78.255 81.100 ;
        RECT 79.020 80.365 79.720 89.860 ;
        RECT 87.845 88.975 88.745 89.935 ;
        RECT 89.285 89.585 90.415 90.755 ;
        RECT 91.000 90.750 91.140 91.435 ;
        RECT 91.635 91.090 92.765 92.260 ;
        RECT 93.160 91.920 94.060 92.330 ;
        RECT 94.500 91.920 94.640 93.040 ;
        RECT 93.160 91.780 94.640 91.920 ;
        RECT 93.160 91.370 94.060 91.780 ;
        RECT 91.000 90.535 91.945 90.750 ;
        RECT 93.540 90.535 93.680 91.370 ;
        RECT 91.000 90.395 93.680 90.535 ;
        RECT 91.000 90.200 91.945 90.395 ;
        RECT 91.045 89.790 91.945 90.200 ;
        RECT 86.070 87.425 87.200 88.595 ;
        RECT 88.225 87.575 88.365 88.975 ;
        RECT 87.845 87.165 88.745 87.575 ;
        RECT 87.805 86.615 88.745 87.165 ;
        RECT 87.805 84.385 87.945 86.615 ;
        RECT 88.605 85.045 89.735 86.215 ;
        RECT 90.180 85.665 91.080 86.110 ;
        RECT 90.180 85.525 92.805 85.665 ;
        RECT 90.180 85.150 91.080 85.525 ;
        RECT 90.325 84.385 90.465 85.150 ;
        RECT 87.805 84.245 90.465 84.385 ;
        RECT 89.820 81.105 89.960 84.245 ;
        RECT 90.680 83.620 91.810 84.790 ;
        RECT 92.665 84.590 92.805 85.525 ;
        RECT 92.285 83.630 93.185 84.590 ;
        RECT 90.680 81.675 91.810 82.845 ;
        RECT 92.490 82.355 93.390 82.765 ;
        RECT 92.405 81.805 93.390 82.355 ;
        RECT 92.405 81.105 92.545 81.805 ;
        RECT 89.820 80.965 92.545 81.105 ;
        RECT 76.920 79.665 79.720 80.365 ;
        RECT 76.920 78.890 77.620 79.665 ;
        RECT 76.850 77.930 77.750 78.890 ;
        RECT 43.900 72.010 45.030 73.180 ;
        RECT 52.885 71.985 54.015 73.155 ;
        RECT 49.725 71.140 50.625 71.160 ;
        RECT 48.995 71.000 50.625 71.140 ;
        RECT 48.995 64.575 49.135 71.000 ;
        RECT 49.725 70.200 50.625 71.000 ;
        RECT 59.480 70.150 60.180 75.385 ;
        RECT 69.525 75.155 70.425 76.115 ;
        RECT 63.380 72.130 64.510 73.300 ;
        RECT 69.625 70.150 70.325 75.155 ;
        RECT 72.020 71.830 73.150 73.000 ;
        RECT 77.510 71.580 78.410 72.540 ;
        RECT 77.675 70.150 78.375 71.580 ;
        RECT 79.020 70.150 79.720 79.665 ;
        RECT 91.470 79.365 91.610 80.965 ;
        RECT 92.950 80.135 94.080 81.305 ;
        RECT 94.570 80.345 95.470 81.305 ;
        RECT 94.950 79.365 95.090 80.345 ;
        RECT 96.105 80.135 97.235 81.305 ;
        RECT 91.470 79.225 95.090 79.365 ;
        RECT 102.215 77.615 102.355 96.010 ;
        RECT 112.445 94.000 112.585 96.010 ;
        RECT 112.900 94.380 114.030 95.550 ;
        RECT 114.830 95.250 114.970 96.010 ;
        RECT 114.470 94.290 115.370 95.250 ;
        RECT 102.700 91.970 103.830 93.140 ;
        RECT 110.995 92.655 112.125 93.825 ;
        RECT 112.445 93.450 113.440 94.000 ;
        RECT 112.540 93.040 113.440 93.450 ;
        RECT 106.555 91.435 109.470 91.575 ;
        RECT 106.555 89.935 106.695 91.435 ;
        RECT 106.175 88.975 107.075 89.935 ;
        RECT 107.615 89.585 108.745 90.755 ;
        RECT 109.330 90.750 109.470 91.435 ;
        RECT 109.965 91.090 111.095 92.260 ;
        RECT 111.490 91.920 112.390 92.330 ;
        RECT 112.830 91.920 112.970 93.040 ;
        RECT 111.490 91.780 112.970 91.920 ;
        RECT 111.490 91.370 112.390 91.780 ;
        RECT 109.330 90.535 110.275 90.750 ;
        RECT 111.870 90.535 112.010 91.370 ;
        RECT 109.330 90.395 112.010 90.535 ;
        RECT 109.330 90.200 110.275 90.395 ;
        RECT 109.375 89.790 110.275 90.200 ;
        RECT 104.400 87.445 105.530 88.615 ;
        RECT 106.555 87.575 106.695 88.975 ;
        RECT 106.175 87.165 107.075 87.575 ;
        RECT 106.135 86.615 107.075 87.165 ;
        RECT 106.135 84.385 106.275 86.615 ;
        RECT 106.935 85.045 108.065 86.215 ;
        RECT 108.510 85.665 109.410 86.110 ;
        RECT 108.510 85.525 111.135 85.665 ;
        RECT 108.510 85.150 109.410 85.525 ;
        RECT 108.655 84.385 108.795 85.150 ;
        RECT 106.135 84.245 108.795 84.385 ;
        RECT 108.150 81.105 108.290 84.245 ;
        RECT 109.010 83.620 110.140 84.790 ;
        RECT 110.995 84.590 111.135 85.525 ;
        RECT 110.615 83.630 111.515 84.590 ;
        RECT 109.010 81.675 110.140 82.845 ;
        RECT 110.820 82.355 111.720 82.765 ;
        RECT 110.735 81.805 111.720 82.355 ;
        RECT 110.735 81.105 110.875 81.805 ;
        RECT 108.150 80.965 110.875 81.105 ;
        RECT 109.800 79.365 109.940 80.965 ;
        RECT 111.280 80.135 112.410 81.305 ;
        RECT 112.900 80.345 113.800 81.305 ;
        RECT 113.280 79.365 113.420 80.345 ;
        RECT 114.435 80.135 115.565 81.305 ;
        RECT 109.800 79.225 113.420 79.365 ;
        RECT 94.040 77.475 114.960 77.615 ;
        RECT 94.040 75.710 94.180 77.475 ;
        RECT 94.330 76.090 95.460 77.260 ;
        RECT 96.055 76.960 96.195 77.475 ;
        RECT 95.850 76.000 96.750 76.960 ;
        RECT 92.375 74.365 93.505 75.535 ;
        RECT 93.920 74.750 94.820 75.710 ;
        RECT 112.475 75.465 112.615 77.475 ;
        RECT 112.930 75.845 114.060 77.015 ;
        RECT 114.820 76.715 114.960 77.475 ;
        RECT 114.500 75.755 115.400 76.715 ;
        RECT 87.935 73.145 90.850 73.285 ;
        RECT 87.935 71.645 88.075 73.145 ;
        RECT 87.555 70.685 88.455 71.645 ;
        RECT 88.995 71.295 90.125 72.465 ;
        RECT 90.710 72.460 90.850 73.145 ;
        RECT 91.345 72.800 92.475 73.970 ;
        RECT 92.870 73.630 93.770 74.040 ;
        RECT 94.210 73.630 94.350 74.750 ;
        RECT 111.025 74.120 112.155 75.290 ;
        RECT 112.475 74.915 113.470 75.465 ;
        RECT 112.570 74.505 113.470 74.915 ;
        RECT 92.870 73.490 94.350 73.630 ;
        RECT 92.870 73.080 93.770 73.490 ;
        RECT 90.710 72.245 91.655 72.460 ;
        RECT 93.250 72.245 93.390 73.080 ;
        RECT 90.710 72.105 93.390 72.245 ;
        RECT 106.585 72.900 109.500 73.040 ;
        RECT 90.710 71.910 91.655 72.105 ;
        RECT 90.755 71.500 91.655 71.910 ;
        RECT 106.585 71.400 106.725 72.900 ;
        RECT 59.480 69.450 79.720 70.150 ;
        RECT 56.375 68.350 57.105 69.120 ;
        RECT 61.105 67.780 61.245 69.450 ;
        RECT 61.720 67.780 62.620 68.190 ;
        RECT 72.480 67.855 73.180 69.450 ;
        RECT 85.780 69.155 86.910 70.325 ;
        RECT 87.935 69.285 88.075 70.685 ;
        RECT 106.205 70.440 107.105 71.400 ;
        RECT 107.645 71.050 108.775 72.220 ;
        RECT 109.360 72.215 109.500 72.900 ;
        RECT 109.995 72.555 111.125 73.725 ;
        RECT 111.520 73.385 112.420 73.795 ;
        RECT 112.860 73.385 113.000 74.505 ;
        RECT 111.520 73.245 113.000 73.385 ;
        RECT 111.520 72.835 112.420 73.245 ;
        RECT 109.360 72.000 110.305 72.215 ;
        RECT 111.900 72.000 112.040 72.835 ;
        RECT 109.360 71.860 112.040 72.000 ;
        RECT 109.360 71.665 110.305 71.860 ;
        RECT 109.405 71.255 110.305 71.665 ;
        RECT 87.555 68.875 88.455 69.285 ;
        RECT 104.430 68.925 105.560 70.095 ;
        RECT 106.585 69.040 106.725 70.440 ;
        RECT 87.515 68.325 88.455 68.875 ;
        RECT 106.205 68.630 107.105 69.040 ;
        RECT 61.105 67.640 62.620 67.780 ;
        RECT 49.495 64.810 50.625 65.980 ;
        RECT 61.105 65.810 61.245 67.640 ;
        RECT 61.720 67.230 62.620 67.640 ;
        RECT 61.720 65.810 62.620 66.370 ;
        RECT 61.105 65.670 62.620 65.810 ;
        RECT 87.515 65.720 87.655 68.325 ;
        RECT 106.165 68.080 107.105 68.630 ;
        RECT 88.315 66.755 89.445 67.925 ;
        RECT 89.890 67.000 90.790 67.820 ;
        RECT 89.890 66.860 92.515 67.000 ;
        RECT 90.035 65.720 90.175 66.860 ;
        RECT 49.725 64.575 50.625 64.620 ;
        RECT 48.995 64.435 50.625 64.575 ;
        RECT 45.935 58.315 46.665 59.085 ;
        RECT 48.995 57.855 49.135 64.435 ;
        RECT 49.725 63.660 50.625 64.435 ;
        RECT 61.105 64.160 61.245 65.670 ;
        RECT 61.720 65.410 62.620 65.670 ;
        RECT 83.440 65.580 90.175 65.720 ;
        RECT 61.720 64.160 62.620 64.550 ;
        RECT 61.105 64.020 62.620 64.160 ;
        RECT 61.105 62.295 61.245 64.020 ;
        RECT 61.720 63.590 62.620 64.020 ;
        RECT 61.730 62.295 62.630 62.735 ;
        RECT 61.105 62.155 62.630 62.295 ;
        RECT 61.105 60.490 61.245 62.155 ;
        RECT 61.730 61.775 62.630 62.155 ;
        RECT 61.730 60.490 62.630 60.910 ;
        RECT 61.105 60.350 62.630 60.490 ;
        RECT 49.495 58.120 50.625 59.290 ;
        RECT 61.105 58.665 61.245 60.350 ;
        RECT 61.730 59.950 62.630 60.350 ;
        RECT 61.730 58.665 62.630 59.085 ;
        RECT 61.105 58.525 62.630 58.665 ;
        RECT 49.725 57.855 50.625 57.925 ;
        RECT 48.995 57.715 50.625 57.855 ;
        RECT 48.995 57.205 49.135 57.715 ;
        RECT 35.590 56.505 49.135 57.205 ;
        RECT 49.725 56.965 50.625 57.715 ;
        RECT 48.995 50.965 49.135 56.505 ;
        RECT 61.105 56.740 61.245 58.525 ;
        RECT 61.730 58.125 62.630 58.525 ;
        RECT 61.720 56.740 62.620 57.275 ;
        RECT 61.105 56.600 62.620 56.740 ;
        RECT 59.425 54.490 60.325 55.450 ;
        RECT 61.105 55.115 61.245 56.600 ;
        RECT 61.720 56.315 62.620 56.600 ;
        RECT 61.730 55.115 62.630 55.450 ;
        RECT 61.105 54.975 62.630 55.115 ;
        RECT 61.730 54.490 62.630 54.975 ;
        RECT 59.805 52.980 59.945 54.490 ;
        RECT 71.145 54.365 71.875 55.135 ;
        RECT 59.805 52.840 62.455 52.980 ;
        RECT 49.495 51.455 50.625 52.625 ;
        RECT 62.315 51.485 62.455 52.840 ;
        RECT 61.955 51.085 62.855 51.485 ;
        RECT 49.650 50.965 50.550 50.995 ;
        RECT 48.995 50.825 50.550 50.965 ;
        RECT 49.650 50.035 50.550 50.825 ;
        RECT 61.340 50.945 62.855 51.085 ;
        RECT 59.510 49.565 60.640 50.735 ;
        RECT 57.995 48.240 59.125 49.410 ;
        RECT 61.340 49.105 61.480 50.945 ;
        RECT 61.955 50.525 62.855 50.945 ;
        RECT 71.145 50.615 71.875 51.385 ;
        RECT 61.955 49.105 62.855 49.665 ;
        RECT 61.340 48.965 62.855 49.105 ;
        RECT 59.510 47.680 60.640 48.850 ;
        RECT 61.340 47.455 61.480 48.965 ;
        RECT 61.955 48.705 62.855 48.965 ;
        RECT 71.045 48.680 72.175 49.850 ;
        RECT 61.955 47.455 62.855 47.845 ;
        RECT 61.340 47.315 62.855 47.455 ;
        RECT 35.530 46.435 36.230 46.485 ;
        RECT 35.530 45.735 42.615 46.435 ;
        RECT 41.915 44.695 42.615 45.735 ;
        RECT 49.495 44.830 50.625 46.000 ;
        RECT 59.510 45.855 60.640 47.025 ;
        RECT 61.340 45.590 61.480 47.315 ;
        RECT 61.955 46.885 62.855 47.315 ;
        RECT 70.985 46.110 72.115 47.280 ;
        RECT 61.965 45.590 62.865 46.025 ;
        RECT 61.340 45.450 62.865 45.590 ;
        RECT 41.815 44.560 42.715 44.695 ;
        RECT 46.390 44.575 47.290 44.690 ;
        RECT 46.390 44.560 54.845 44.575 ;
        RECT 41.815 43.875 54.845 44.560 ;
        RECT 59.510 43.980 60.640 45.150 ;
        RECT 41.815 43.860 47.290 43.875 ;
        RECT 41.815 43.735 42.715 43.860 ;
        RECT 37.420 38.600 38.550 39.770 ;
        RECT 41.835 37.705 42.735 38.035 ;
        RECT 42.945 37.705 43.085 43.860 ;
        RECT 41.835 37.405 43.085 37.705 ;
        RECT 41.835 37.075 42.735 37.405 ;
        RECT 37.070 31.895 38.200 33.065 ;
        RECT 41.795 31.385 42.695 31.920 ;
        RECT 42.945 31.385 43.085 37.405 ;
        RECT 41.795 31.085 43.085 31.385 ;
        RECT 41.795 30.960 42.695 31.085 ;
        RECT 21.320 27.400 23.690 29.730 ;
        RECT 37.070 25.780 38.200 26.950 ;
        RECT 41.835 24.895 42.735 25.495 ;
        RECT 42.945 24.895 43.085 31.085 ;
        RECT 41.835 24.755 43.085 24.895 ;
        RECT 44.390 42.220 44.690 43.860 ;
        RECT 46.390 43.730 47.290 43.860 ;
        RECT 44.890 42.220 45.790 42.550 ;
        RECT 44.390 41.920 45.790 42.220 ;
        RECT 44.390 37.730 44.690 41.920 ;
        RECT 44.890 41.590 45.790 41.920 ;
        RECT 46.230 38.610 47.360 39.780 ;
        RECT 46.390 37.730 47.290 38.060 ;
        RECT 44.390 37.430 47.290 37.730 ;
        RECT 44.390 35.255 44.690 37.430 ;
        RECT 46.390 37.100 47.290 37.430 ;
        RECT 54.145 35.865 54.845 43.875 ;
        RECT 61.340 43.785 61.480 45.450 ;
        RECT 61.965 45.065 62.865 45.450 ;
        RECT 61.965 43.785 62.865 44.205 ;
        RECT 61.340 43.645 62.865 43.785 ;
        RECT 59.510 42.160 60.640 43.330 ;
        RECT 61.340 41.960 61.480 43.645 ;
        RECT 61.965 43.245 62.865 43.645 ;
        RECT 71.095 43.605 72.225 44.775 ;
        RECT 61.965 41.960 62.865 42.380 ;
        RECT 61.340 41.820 62.865 41.960 ;
        RECT 59.510 40.420 60.640 41.590 ;
        RECT 61.340 40.155 61.480 41.820 ;
        RECT 61.965 41.420 62.865 41.820 ;
        RECT 71.095 40.995 72.225 42.165 ;
        RECT 61.955 40.155 62.855 40.570 ;
        RECT 61.340 40.015 62.855 40.155 ;
        RECT 59.510 38.585 60.640 39.755 ;
        RECT 61.340 38.335 61.480 40.015 ;
        RECT 61.955 39.610 62.855 40.015 ;
        RECT 61.965 38.335 62.865 38.745 ;
        RECT 71.095 38.510 72.225 39.680 ;
        RECT 61.340 38.195 62.865 38.335 ;
        RECT 61.965 37.785 62.865 38.195 ;
        RECT 71.180 37.025 71.910 37.795 ;
        RECT 83.440 37.275 83.580 65.580 ;
        RECT 89.700 62.865 89.840 65.580 ;
        RECT 90.390 65.330 91.520 66.500 ;
        RECT 92.375 66.300 92.515 66.860 ;
        RECT 91.995 65.340 92.895 66.300 ;
        RECT 106.165 65.850 106.305 68.080 ;
        RECT 106.965 66.510 108.095 67.680 ;
        RECT 108.540 67.130 109.440 67.575 ;
        RECT 108.540 66.990 111.165 67.130 ;
        RECT 108.540 66.615 109.440 66.990 ;
        RECT 108.685 65.850 108.825 66.615 ;
        RECT 106.165 65.710 108.825 65.850 ;
        RECT 90.390 63.385 91.520 64.555 ;
        RECT 92.200 64.065 93.100 64.475 ;
        RECT 91.910 63.925 93.100 64.065 ;
        RECT 91.910 62.865 92.050 63.925 ;
        RECT 92.200 63.515 93.100 63.925 ;
        RECT 89.700 62.725 92.050 62.865 ;
        RECT 91.180 60.700 91.320 62.725 ;
        RECT 92.660 61.845 93.790 63.015 ;
        RECT 94.280 62.055 95.180 63.015 ;
        RECT 94.660 60.700 94.800 62.055 ;
        RECT 95.815 61.845 96.945 63.015 ;
        RECT 108.180 62.570 108.320 65.710 ;
        RECT 109.040 65.085 110.170 66.255 ;
        RECT 111.025 66.055 111.165 66.990 ;
        RECT 110.645 65.095 111.545 66.055 ;
        RECT 109.040 63.140 110.170 64.310 ;
        RECT 110.850 63.820 111.750 64.230 ;
        RECT 110.765 63.270 111.750 63.820 ;
        RECT 110.765 62.570 110.905 63.270 ;
        RECT 108.180 62.430 110.905 62.570 ;
        RECT 91.180 60.560 94.800 60.700 ;
        RECT 109.830 60.830 109.970 62.430 ;
        RECT 111.310 61.600 112.440 62.770 ;
        RECT 112.930 61.810 113.830 62.770 ;
        RECT 113.310 60.830 113.450 61.810 ;
        RECT 114.465 61.600 115.595 62.770 ;
        RECT 109.830 60.690 113.450 60.830 ;
        RECT 94.660 60.465 94.800 60.560 ;
        RECT 94.660 60.325 94.840 60.465 ;
        RECT 94.700 59.410 94.840 60.325 ;
        RECT 94.700 59.270 101.780 59.410 ;
        RECT 101.640 39.370 101.780 59.270 ;
        RECT 105.295 57.670 112.970 58.370 ;
        RECT 105.295 57.140 105.995 57.670 ;
        RECT 108.325 57.140 109.025 57.670 ;
        RECT 112.270 57.140 112.970 57.670 ;
        RECT 105.195 57.010 106.095 57.140 ;
        RECT 102.765 56.310 106.095 57.010 ;
        RECT 102.765 51.760 103.465 56.310 ;
        RECT 105.195 56.180 106.095 56.310 ;
        RECT 106.665 55.965 107.795 57.135 ;
        RECT 108.200 56.180 109.100 57.140 ;
        RECT 109.665 55.965 110.795 57.135 ;
        RECT 112.170 56.180 113.070 57.140 ;
        RECT 104.415 54.555 105.545 55.725 ;
        RECT 104.080 52.880 105.210 54.050 ;
        RECT 105.750 53.105 106.650 54.065 ;
        RECT 105.950 52.085 106.650 53.105 ;
        RECT 104.810 51.890 106.650 52.085 ;
        RECT 104.710 51.760 106.650 51.890 ;
        RECT 102.705 51.385 106.650 51.760 ;
        RECT 102.705 51.060 105.610 51.385 ;
        RECT 102.705 48.480 103.405 51.060 ;
        RECT 104.710 50.930 105.610 51.060 ;
        RECT 104.080 49.260 105.210 50.430 ;
        RECT 104.710 48.480 105.610 48.610 ;
        RECT 102.705 48.275 105.610 48.480 ;
        RECT 102.690 47.780 105.610 48.275 ;
        RECT 102.690 47.575 103.405 47.780 ;
        RECT 104.710 47.650 105.610 47.780 ;
        RECT 102.690 41.950 103.390 47.575 ;
        RECT 104.080 45.510 105.210 46.680 ;
        RECT 105.750 45.610 106.650 46.570 ;
        RECT 104.755 43.905 105.885 45.075 ;
        RECT 106.130 43.440 106.270 45.610 ;
        RECT 105.750 42.480 106.650 43.440 ;
        RECT 106.115 41.950 106.255 42.480 ;
        RECT 107.165 42.415 108.295 43.585 ;
        RECT 108.650 42.455 109.550 43.415 ;
        RECT 109.895 42.455 111.025 43.625 ;
        RECT 112.170 43.490 113.070 43.670 ;
        RECT 112.170 43.440 123.875 43.490 ;
        RECT 112.170 42.800 124.100 43.440 ;
        RECT 112.170 42.790 123.875 42.800 ;
        RECT 112.170 42.710 113.070 42.790 ;
        RECT 102.690 41.705 106.605 41.950 ;
        RECT 108.715 41.705 109.415 42.455 ;
        RECT 112.270 41.705 112.970 42.710 ;
        RECT 102.690 41.250 112.970 41.705 ;
        RECT 106.185 41.005 112.970 41.250 ;
        RECT 110.830 39.370 111.430 39.620 ;
        RECT 101.640 39.230 111.430 39.370 ;
        RECT 110.830 38.980 111.430 39.230 ;
        RECT 83.420 37.135 83.580 37.275 ;
        RECT 56.165 36.275 69.730 36.975 ;
        RECT 56.165 35.995 56.865 36.275 ;
        RECT 55.850 35.865 56.865 35.995 ;
        RECT 44.890 35.255 45.790 35.585 ;
        RECT 44.390 34.955 45.790 35.255 ;
        RECT 54.145 35.165 56.865 35.865 ;
        RECT 55.850 35.035 56.750 35.165 ;
        RECT 44.390 31.210 44.690 34.955 ;
        RECT 44.890 34.625 45.790 34.955 ;
        RECT 57.070 34.375 58.200 35.545 ;
        RECT 69.030 34.080 69.730 36.275 ;
        RECT 72.485 36.155 73.065 36.350 ;
        RECT 83.420 36.155 83.560 37.135 ;
        RECT 72.485 36.015 83.560 36.155 ;
        RECT 70.910 34.735 72.040 35.905 ;
        RECT 72.485 35.710 73.065 36.015 ;
        RECT 68.930 33.120 69.830 34.080 ;
        RECT 46.215 31.905 47.345 33.075 ;
        RECT 47.580 31.210 48.480 31.900 ;
        RECT 57.070 31.330 58.200 32.500 ;
        RECT 44.390 31.070 48.480 31.210 ;
        RECT 44.390 28.970 44.690 31.070 ;
        RECT 47.580 30.940 48.480 31.070 ;
        RECT 44.890 28.970 45.790 29.300 ;
        RECT 44.390 28.670 45.790 28.970 ;
        RECT 44.390 25.100 44.690 28.670 ;
        RECT 44.890 28.340 45.790 28.670 ;
        RECT 46.250 25.810 47.380 26.980 ;
        RECT 47.580 25.100 48.480 25.495 ;
        RECT 44.390 24.800 48.480 25.100 ;
        RECT 41.835 24.535 42.735 24.755 ;
        RECT 45.190 23.225 45.490 24.800 ;
        RECT 47.580 24.535 48.480 24.800 ;
        RECT 44.890 22.265 45.790 23.225 ;
        RECT 36.080 19.385 37.210 20.555 ;
        RECT 46.205 19.405 47.335 20.575 ;
        RECT 95.290 17.535 96.420 18.705 ;
        RECT 138.170 14.665 140.540 16.995 ;
        RECT 138.570 8.825 140.140 10.355 ;
        RECT 128.240 6.615 129.810 8.145 ;
        RECT 106.305 4.695 107.875 6.225 ;
        RECT 83.965 3.030 85.535 4.560 ;
        RECT 61.790 1.490 63.360 3.020 ;
      LAYER met3 ;
        RECT 97.740 213.665 98.040 213.670 ;
        RECT 97.525 212.895 98.255 213.665 ;
        RECT 105.720 213.035 106.450 213.805 ;
        RECT 97.740 209.495 98.040 212.895 ;
        RECT 105.935 209.495 106.235 213.035 ;
        RECT 97.740 209.195 106.235 209.495 ;
        RECT 97.740 206.490 98.040 209.195 ;
        RECT 105.935 206.725 106.235 209.195 ;
        RECT 97.525 205.720 98.255 206.490 ;
        RECT 105.720 205.955 106.450 206.725 ;
        RECT 97.740 199.540 98.040 205.720 ;
        RECT 105.935 199.855 106.235 205.955 ;
        RECT 97.525 198.770 98.255 199.540 ;
        RECT 105.720 199.085 106.450 199.855 ;
        RECT 97.740 192.515 98.040 198.770 ;
        RECT 105.935 192.515 106.235 199.085 ;
        RECT 95.755 192.230 96.485 192.465 ;
        RECT 97.525 192.230 98.255 192.515 ;
        RECT 95.755 191.930 98.255 192.230 ;
        RECT 95.755 191.695 96.485 191.930 ;
        RECT 97.525 191.745 98.255 191.930 ;
        RECT 105.720 191.745 106.450 192.515 ;
        RECT 53.170 190.085 54.300 190.585 ;
        RECT 53.170 189.785 57.445 190.085 ;
        RECT 53.170 189.415 54.300 189.785 ;
        RECT 57.145 188.285 57.445 189.785 ;
        RECT 97.525 188.715 98.255 189.485 ;
        RECT 97.740 188.285 98.040 188.715 ;
        RECT 57.145 187.985 98.040 188.285 ;
        RECT 105.935 173.450 106.235 191.745 ;
        RECT 105.690 172.680 106.420 173.450 ;
        RECT 105.935 166.660 106.235 172.680 ;
        RECT 105.690 165.890 106.420 166.660 ;
        RECT 17.610 148.645 19.990 148.805 ;
        RECT 21.320 148.645 23.690 148.810 ;
        RECT 17.610 146.645 23.690 148.645 ;
        RECT 17.610 146.485 19.990 146.645 ;
        RECT 21.320 146.480 23.690 146.645 ;
        RECT 138.170 147.660 140.540 147.825 ;
        RECT 143.700 147.660 146.080 147.820 ;
        RECT 138.170 145.660 146.080 147.660 ;
        RECT 138.170 145.495 140.540 145.660 ;
        RECT 143.700 145.500 146.080 145.660 ;
        RECT 71.590 108.720 72.320 108.840 ;
        RECT 42.230 108.705 72.320 108.720 ;
        RECT 40.880 108.420 72.320 108.705 ;
        RECT 40.880 108.405 42.530 108.420 ;
        RECT 40.880 101.500 41.180 108.405 ;
        RECT 71.590 108.070 72.320 108.420 ;
        RECT 43.900 101.500 45.030 102.250 ;
        RECT 40.880 101.200 45.030 101.500 ;
        RECT 40.880 91.630 41.180 101.200 ;
        RECT 43.900 101.080 45.030 101.200 ;
        RECT 52.885 101.115 54.015 102.285 ;
        RECT 53.300 99.610 53.600 101.115 ;
        RECT 63.380 101.055 64.510 102.225 ;
        RECT 63.565 100.035 63.865 101.055 ;
        RECT 51.635 99.310 53.600 99.610 ;
        RECT 62.000 99.735 63.945 100.035 ;
        RECT 43.900 91.630 45.030 92.340 ;
        RECT 40.880 91.330 45.030 91.630 ;
        RECT 43.900 91.170 45.030 91.330 ;
        RECT 51.635 92.050 51.935 99.310 ;
        RECT 52.885 92.050 54.015 92.375 ;
        RECT 51.635 91.750 54.015 92.050 ;
        RECT 43.900 81.535 45.030 82.185 ;
        RECT 42.935 81.235 45.030 81.535 ;
        RECT 42.935 72.625 43.235 81.235 ;
        RECT 43.900 81.015 45.030 81.235 ;
        RECT 51.635 81.925 51.935 91.750 ;
        RECT 52.885 91.205 54.015 91.750 ;
        RECT 62.000 91.770 62.300 99.735 ;
        RECT 120.125 97.885 120.855 97.920 ;
        RECT 102.875 97.185 120.855 97.885 ;
        RECT 94.570 95.355 95.700 95.550 ;
        RECT 92.880 94.655 95.700 95.355 ;
        RECT 92.880 93.825 93.580 94.655 ;
        RECT 94.570 94.380 95.700 94.655 ;
        RECT 92.665 93.600 93.795 93.825 ;
        RECT 91.545 92.900 93.795 93.600 ;
        RECT 102.875 93.140 103.575 97.185 ;
        RECT 120.125 97.150 120.855 97.185 ;
        RECT 112.900 95.355 114.030 95.550 ;
        RECT 111.210 94.655 114.030 95.355 ;
        RECT 111.210 93.825 111.910 94.655 ;
        RECT 112.900 94.380 114.030 94.655 ;
        RECT 110.995 93.600 112.125 93.825 ;
        RECT 63.380 91.770 64.510 92.330 ;
        RECT 91.545 92.260 92.245 92.900 ;
        RECT 92.665 92.655 93.795 92.900 ;
        RECT 91.545 92.245 92.765 92.260 ;
        RECT 62.000 91.470 64.510 91.770 ;
        RECT 52.885 81.925 54.015 82.360 ;
        RECT 51.635 81.625 54.015 81.925 ;
        RECT 50.455 75.780 51.185 76.015 ;
        RECT 51.635 75.780 51.935 81.625 ;
        RECT 52.885 81.190 54.015 81.625 ;
        RECT 62.000 82.020 62.300 91.470 ;
        RECT 63.380 91.160 64.510 91.470 ;
        RECT 89.500 91.545 92.765 92.245 ;
        RECT 102.700 91.970 103.830 93.140 ;
        RECT 109.960 92.900 112.125 93.600 ;
        RECT 109.960 92.330 110.660 92.900 ;
        RECT 110.995 92.655 112.125 92.900 ;
        RECT 107.830 92.260 110.880 92.330 ;
        RECT 89.500 90.755 90.200 91.545 ;
        RECT 91.635 91.090 92.765 91.545 ;
        RECT 107.830 91.630 111.095 92.260 ;
        RECT 107.830 90.755 108.530 91.630 ;
        RECT 109.965 91.090 111.095 91.630 ;
        RECT 89.285 90.375 90.415 90.755 ;
        RECT 107.615 90.460 108.745 90.755 ;
        RECT 86.330 89.675 90.415 90.375 ;
        RECT 86.330 88.595 87.030 89.675 ;
        RECT 89.285 89.585 90.415 89.675 ;
        RECT 104.660 89.760 108.745 90.460 ;
        RECT 104.660 88.615 105.360 89.760 ;
        RECT 107.615 89.585 108.745 89.760 ;
        RECT 86.070 87.425 87.200 88.595 ;
        RECT 104.400 87.445 105.530 88.615 ;
        RECT 86.345 85.840 87.045 87.425 ;
        RECT 88.605 85.840 89.735 86.215 ;
        RECT 86.345 85.140 89.735 85.840 ;
        RECT 104.675 85.980 105.375 87.445 ;
        RECT 106.935 85.980 108.065 86.215 ;
        RECT 104.675 85.280 108.065 85.980 ;
        RECT 88.605 85.045 89.735 85.140 ;
        RECT 106.935 85.045 108.065 85.280 ;
        RECT 88.960 84.065 89.660 85.045 ;
        RECT 90.680 84.065 91.810 84.790 ;
        RECT 88.960 83.620 91.810 84.065 ;
        RECT 107.290 84.205 107.990 85.045 ;
        RECT 109.010 84.205 110.140 84.790 ;
        RECT 107.290 83.620 110.140 84.205 ;
        RECT 88.960 83.365 91.595 83.620 ;
        RECT 107.290 83.505 109.925 83.620 ;
        RECT 90.895 82.845 91.595 83.365 ;
        RECT 109.225 82.845 109.925 83.505 ;
        RECT 63.380 82.020 64.510 82.475 ;
        RECT 72.425 82.225 73.555 82.625 ;
        RECT 62.000 81.720 64.510 82.020 ;
        RECT 50.455 75.480 51.935 75.780 ;
        RECT 50.455 75.245 51.185 75.480 ;
        RECT 43.900 72.745 45.030 73.180 ;
        RECT 51.635 73.045 51.935 75.480 ;
        RECT 52.885 73.055 54.015 73.155 ;
        RECT 62.000 73.055 62.300 81.720 ;
        RECT 63.380 81.305 64.510 81.720 ;
        RECT 70.875 81.925 73.555 82.225 ;
        RECT 63.380 73.055 64.510 73.300 ;
        RECT 52.885 73.045 64.510 73.055 ;
        RECT 51.635 72.755 64.510 73.045 ;
        RECT 51.635 72.745 54.015 72.755 ;
        RECT 43.900 72.625 51.935 72.745 ;
        RECT 42.935 72.445 51.935 72.625 ;
        RECT 42.935 72.325 45.030 72.445 ;
        RECT 43.900 72.010 45.030 72.325 ;
        RECT 52.885 71.985 54.015 72.745 ;
        RECT 63.380 72.130 64.510 72.755 ;
        RECT 70.875 72.535 71.175 81.925 ;
        RECT 72.425 81.455 73.555 81.925 ;
        RECT 90.680 81.675 91.810 82.845 ;
        RECT 109.010 81.675 110.140 82.845 ;
        RECT 90.760 80.930 91.460 81.675 ;
        RECT 92.950 80.930 94.080 81.305 ;
        RECT 90.760 80.230 94.080 80.930 ;
        RECT 92.950 80.135 94.080 80.230 ;
        RECT 96.105 80.950 97.235 81.305 ;
        RECT 109.090 80.950 109.790 81.675 ;
        RECT 111.280 80.950 112.410 81.305 ;
        RECT 96.105 80.250 112.410 80.950 ;
        RECT 96.105 80.135 97.235 80.250 ;
        RECT 93.165 79.810 93.865 80.135 ;
        RECT 96.330 79.810 97.030 80.135 ;
        RECT 93.165 79.110 97.030 79.810 ;
        RECT 94.330 77.065 95.460 77.260 ;
        RECT 92.590 76.365 95.460 77.065 ;
        RECT 92.590 75.535 93.290 76.365 ;
        RECT 94.330 76.090 95.460 76.365 ;
        RECT 92.375 75.310 93.505 75.535 ;
        RECT 91.360 74.610 93.505 75.310 ;
        RECT 91.360 74.100 92.060 74.610 ;
        RECT 92.375 74.365 93.505 74.610 ;
        RECT 89.015 73.970 92.065 74.100 ;
        RECT 89.015 73.400 92.475 73.970 ;
        RECT 72.020 72.535 73.150 73.000 ;
        RECT 70.875 72.235 73.150 72.535 ;
        RECT 89.015 72.465 89.715 73.400 ;
        RECT 91.345 72.800 92.475 73.400 ;
        RECT 70.875 71.685 71.175 72.235 ;
        RECT 72.020 71.830 73.150 72.235 ;
        RECT 88.995 72.230 90.125 72.465 ;
        RECT 48.605 71.385 71.175 71.685 ;
        RECT 85.845 71.530 90.125 72.230 ;
        RECT 48.605 65.545 48.905 71.385 ;
        RECT 56.560 69.120 56.860 71.385 ;
        RECT 85.845 70.325 86.545 71.530 ;
        RECT 88.995 71.295 90.125 71.530 ;
        RECT 85.780 69.155 86.910 70.325 ;
        RECT 56.375 68.350 57.105 69.120 ;
        RECT 85.845 67.460 86.545 69.155 ;
        RECT 88.315 67.460 89.445 67.925 ;
        RECT 85.845 66.760 89.445 67.460 ;
        RECT 88.315 66.755 89.445 66.760 ;
        RECT 49.495 65.545 50.625 65.980 ;
        RECT 48.605 65.245 50.625 65.545 ;
        RECT 45.935 58.805 46.665 59.085 ;
        RECT 48.605 58.805 48.905 65.245 ;
        RECT 49.495 64.810 50.625 65.245 ;
        RECT 88.670 65.685 89.370 66.755 ;
        RECT 90.390 65.685 91.520 66.500 ;
        RECT 88.670 65.330 91.520 65.685 ;
        RECT 88.670 64.985 91.305 65.330 ;
        RECT 90.605 64.555 91.305 64.985 ;
        RECT 90.390 63.385 91.520 64.555 ;
        RECT 90.470 62.550 91.170 63.385 ;
        RECT 92.660 62.550 93.790 63.015 ;
        RECT 90.470 61.850 93.790 62.550 ;
        RECT 92.660 61.845 93.790 61.850 ;
        RECT 95.815 62.315 96.945 63.015 ;
        RECT 101.435 62.315 102.135 80.250 ;
        RECT 111.280 80.135 112.410 80.250 ;
        RECT 114.435 80.135 115.565 81.305 ;
        RECT 111.625 79.830 112.325 80.135 ;
        RECT 114.650 79.830 115.350 80.135 ;
        RECT 111.625 79.130 115.350 79.830 ;
        RECT 112.930 76.820 114.060 77.015 ;
        RECT 111.240 76.120 114.060 76.820 ;
        RECT 111.240 75.290 111.940 76.120 ;
        RECT 112.930 75.845 114.060 76.120 ;
        RECT 111.025 75.065 112.155 75.290 ;
        RECT 109.985 74.365 112.155 75.065 ;
        RECT 109.985 73.855 110.685 74.365 ;
        RECT 111.025 74.120 112.155 74.365 ;
        RECT 107.645 73.725 110.695 73.855 ;
        RECT 107.645 73.155 111.125 73.725 ;
        RECT 107.645 72.220 108.345 73.155 ;
        RECT 109.985 73.140 111.125 73.155 ;
        RECT 109.995 72.555 111.125 73.140 ;
        RECT 107.645 71.985 108.775 72.220 ;
        RECT 104.475 71.285 108.775 71.985 ;
        RECT 104.475 70.095 105.175 71.285 ;
        RECT 107.645 71.050 108.775 71.285 ;
        RECT 104.430 68.925 105.560 70.095 ;
        RECT 104.475 67.445 105.175 68.925 ;
        RECT 106.965 67.445 108.095 67.680 ;
        RECT 104.475 66.745 108.095 67.445 ;
        RECT 106.965 66.510 108.095 66.745 ;
        RECT 107.320 65.670 108.020 66.510 ;
        RECT 109.040 65.670 110.170 66.255 ;
        RECT 107.320 65.085 110.170 65.670 ;
        RECT 107.320 64.970 109.955 65.085 ;
        RECT 109.255 64.310 109.955 64.970 ;
        RECT 109.040 63.140 110.170 64.310 ;
        RECT 109.120 62.315 109.820 63.140 ;
        RECT 111.310 62.315 112.440 62.770 ;
        RECT 95.815 61.845 112.440 62.315 ;
        RECT 92.875 61.430 93.575 61.845 ;
        RECT 96.030 61.615 112.440 61.845 ;
        RECT 96.030 61.430 96.740 61.615 ;
        RECT 92.875 60.730 96.740 61.430 ;
        RECT 100.545 60.950 101.245 61.615 ;
        RECT 111.310 61.600 112.440 61.615 ;
        RECT 114.465 61.600 115.595 62.770 ;
        RECT 111.525 61.195 112.225 61.600 ;
        RECT 114.690 61.195 115.390 61.600 ;
        RECT 100.545 60.210 101.320 60.950 ;
        RECT 111.525 60.495 115.390 61.195 ;
        RECT 100.600 60.170 101.320 60.210 ;
        RECT 49.495 58.805 50.625 59.290 ;
        RECT 45.935 58.505 50.625 58.805 ;
        RECT 45.935 58.315 46.665 58.505 ;
        RECT 49.495 58.120 50.625 58.505 ;
        RECT 103.310 58.920 107.980 58.950 ;
        RECT 103.310 58.250 110.580 58.920 ;
        RECT 103.310 55.505 104.010 58.250 ;
        RECT 106.900 58.220 110.580 58.250 ;
        RECT 106.900 57.135 107.600 58.220 ;
        RECT 109.880 57.135 110.580 58.220 ;
        RECT 106.665 55.965 107.795 57.135 ;
        RECT 109.665 55.965 110.795 57.135 ;
        RECT 104.415 55.505 105.545 55.725 ;
        RECT 70.950 54.160 72.070 55.340 ;
        RECT 102.115 54.805 105.545 55.505 ;
        RECT 102.115 53.615 102.815 54.805 ;
        RECT 104.415 54.555 105.545 54.805 ;
        RECT 104.080 53.615 105.210 54.050 ;
        RECT 102.115 53.315 105.210 53.615 ;
        RECT 49.495 52.190 50.625 52.625 ;
        RECT 48.595 51.890 50.625 52.190 ;
        RECT 48.595 45.710 48.895 51.890 ;
        RECT 49.495 51.455 50.625 51.890 ;
        RECT 59.510 49.565 60.640 50.735 ;
        RECT 70.950 50.410 72.070 51.590 ;
        RECT 102.115 50.575 102.815 53.315 ;
        RECT 104.080 52.880 105.210 53.315 ;
        RECT 102.115 49.995 102.880 50.575 ;
        RECT 104.080 49.995 105.210 50.430 ;
        RECT 102.115 49.875 105.210 49.995 ;
        RECT 57.995 48.240 59.125 49.410 ;
        RECT 59.925 48.850 60.225 49.565 ;
        RECT 58.535 46.695 58.835 48.240 ;
        RECT 59.510 47.680 60.640 48.850 ;
        RECT 71.045 48.680 72.175 49.850 ;
        RECT 102.175 49.695 105.210 49.875 ;
        RECT 59.925 47.025 60.225 47.680 ;
        RECT 71.510 47.280 71.810 48.680 ;
        RECT 59.510 46.695 60.640 47.025 ;
        RECT 58.535 46.395 60.640 46.695 ;
        RECT 49.495 45.800 50.625 46.000 ;
        RECT 58.535 45.800 58.835 46.395 ;
        RECT 59.510 45.855 60.640 46.395 ;
        RECT 70.985 46.110 72.115 47.280 ;
        RECT 49.495 45.710 58.835 45.800 ;
        RECT 48.595 45.500 58.835 45.710 ;
        RECT 48.595 45.410 50.625 45.500 ;
        RECT 49.495 44.830 50.625 45.410 ;
        RECT 59.925 45.150 60.225 45.855 ;
        RECT 59.510 43.980 60.640 45.150 ;
        RECT 71.510 44.775 71.810 46.110 ;
        RECT 102.175 44.840 102.875 49.695 ;
        RECT 104.080 49.260 105.210 49.695 ;
        RECT 104.080 46.445 105.210 46.680 ;
        RECT 103.735 45.510 105.210 46.445 ;
        RECT 103.735 44.840 104.435 45.510 ;
        RECT 104.755 44.840 105.885 45.075 ;
        RECT 59.925 43.330 60.225 43.980 ;
        RECT 71.095 43.605 72.225 44.775 ;
        RECT 102.175 44.140 105.885 44.840 ;
        RECT 59.510 42.160 60.640 43.330 ;
        RECT 71.510 42.165 71.810 43.605 ;
        RECT 59.925 41.590 60.225 42.160 ;
        RECT 59.510 40.420 60.640 41.590 ;
        RECT 71.095 40.995 72.225 42.165 ;
        RECT 103.735 41.755 104.435 44.140 ;
        RECT 104.755 43.905 105.885 44.140 ;
        RECT 107.165 42.415 108.295 43.585 ;
        RECT 109.895 42.455 111.025 43.625 ;
        RECT 103.735 41.455 104.575 41.755 ;
        RECT 35.030 39.335 36.670 39.365 ;
        RECT 37.420 39.335 38.550 39.770 ;
        RECT 46.230 39.345 47.360 39.780 ;
        RECT 59.925 39.755 60.225 40.420 ;
        RECT 35.030 39.035 38.550 39.335 ;
        RECT 35.030 32.865 35.330 39.035 ;
        RECT 37.420 38.600 38.550 39.035 ;
        RECT 44.055 39.045 47.360 39.345 ;
        RECT 37.070 32.865 38.200 33.065 ;
        RECT 35.030 32.565 38.200 32.865 ;
        RECT 17.610 29.565 19.990 29.725 ;
        RECT 21.320 29.565 23.690 29.730 ;
        RECT 17.610 27.565 23.690 29.565 ;
        RECT 17.610 27.405 19.990 27.565 ;
        RECT 21.320 27.400 23.690 27.565 ;
        RECT 35.030 26.645 35.330 32.565 ;
        RECT 37.070 31.895 38.200 32.565 ;
        RECT 44.055 32.650 44.355 39.045 ;
        RECT 46.230 38.610 47.360 39.045 ;
        RECT 59.510 38.585 60.640 39.755 ;
        RECT 71.510 39.680 71.810 40.995 ;
        RECT 104.075 40.865 104.375 41.455 ;
        RECT 107.380 40.865 108.080 42.415 ;
        RECT 110.095 40.865 110.795 42.455 ;
        RECT 95.400 40.165 110.795 40.865 ;
        RECT 71.095 38.510 72.225 39.680 ;
        RECT 71.510 37.795 71.810 38.510 ;
        RECT 71.180 37.025 71.910 37.795 ;
        RECT 57.070 35.110 58.200 35.545 ;
        RECT 70.910 35.110 72.040 35.905 ;
        RECT 54.255 34.810 72.040 35.110 ;
        RECT 46.215 32.705 47.345 33.075 ;
        RECT 54.255 32.705 54.555 34.810 ;
        RECT 57.070 34.375 58.200 34.810 ;
        RECT 70.910 34.735 72.040 34.810 ;
        RECT 44.055 32.640 45.240 32.650 ;
        RECT 46.215 32.640 54.555 32.705 ;
        RECT 44.055 32.405 54.555 32.640 ;
        RECT 44.055 32.340 47.345 32.405 ;
        RECT 37.070 26.645 38.200 26.950 ;
        RECT 35.030 26.345 38.200 26.645 ;
        RECT 35.030 20.120 35.330 26.345 ;
        RECT 37.070 25.780 38.200 26.345 ;
        RECT 44.055 26.615 44.355 32.340 ;
        RECT 46.215 31.905 47.345 32.340 ;
        RECT 55.885 32.065 56.605 32.190 ;
        RECT 57.070 32.065 58.200 32.500 ;
        RECT 55.885 31.765 58.200 32.065 ;
        RECT 55.885 31.410 56.605 31.765 ;
        RECT 57.070 31.330 58.200 31.765 ;
        RECT 46.250 26.615 47.380 26.980 ;
        RECT 44.055 26.315 47.380 26.615 ;
        RECT 36.080 20.120 37.210 20.555 ;
        RECT 35.030 20.035 37.210 20.120 ;
        RECT 44.055 20.035 44.355 26.315 ;
        RECT 44.985 26.295 45.285 26.315 ;
        RECT 46.250 25.810 47.380 26.315 ;
        RECT 46.205 20.035 47.335 20.575 ;
        RECT 35.030 19.820 47.335 20.035 ;
        RECT 36.080 19.735 47.335 19.820 ;
        RECT 36.080 19.385 37.210 19.735 ;
        RECT 46.205 19.405 47.335 19.735 ;
        RECT 95.400 18.705 96.100 40.165 ;
        RECT 95.290 18.470 96.420 18.705 ;
        RECT 100.090 18.470 122.545 34.770 ;
        RECT 95.290 17.770 122.545 18.470 ;
        RECT 95.290 17.535 96.420 17.770 ;
        RECT 100.090 12.320 122.545 17.770 ;
        RECT 138.170 16.830 140.540 16.995 ;
        RECT 143.700 16.830 146.080 16.990 ;
        RECT 138.170 14.830 146.080 16.830 ;
        RECT 138.170 14.665 140.540 14.830 ;
        RECT 143.700 14.670 146.080 14.830 ;
        RECT 139.355 10.355 144.930 10.590 ;
        RECT 138.570 10.350 144.930 10.355 ;
        RECT 138.570 8.830 145.680 10.350 ;
        RECT 138.570 8.825 144.930 8.830 ;
        RECT 139.355 8.590 144.930 8.825 ;
        RECT 128.240 8.140 134.600 8.380 ;
        RECT 128.240 6.620 135.350 8.140 ;
        RECT 106.305 6.220 112.665 6.460 ;
        RECT 128.240 6.380 134.600 6.620 ;
        RECT 83.965 4.555 90.325 4.795 ;
        RECT 106.305 4.700 113.415 6.220 ;
        RECT 67.320 3.030 68.900 3.050 ;
        RECT 61.790 2.030 68.900 3.030 ;
        RECT 83.965 3.035 91.075 4.555 ;
        RECT 106.305 4.460 112.665 4.700 ;
        RECT 83.965 2.795 90.325 3.035 ;
        RECT 61.790 1.490 63.360 2.030 ;
        RECT 67.320 1.530 68.900 2.030 ;
      LAYER met4 ;
        RECT 3.980 225.065 3.990 225.760 ;
        RECT 7.660 225.065 7.670 225.760 ;
        RECT 11.340 225.065 11.350 225.760 ;
        RECT 15.020 225.065 15.030 225.760 ;
        RECT 18.700 225.065 18.710 225.760 ;
        RECT 22.380 225.065 22.390 225.760 ;
        RECT 26.060 225.065 26.070 225.760 ;
        RECT 29.740 225.065 29.750 225.760 ;
        RECT 33.420 225.065 33.430 225.760 ;
        RECT 37.100 225.065 37.110 225.760 ;
        RECT 40.780 225.065 40.790 225.760 ;
        RECT 44.460 225.065 44.470 225.760 ;
        RECT 48.140 225.065 48.150 225.760 ;
        RECT 51.820 225.065 51.830 225.760 ;
        RECT 55.500 225.065 55.510 225.760 ;
        RECT 59.180 225.065 59.190 225.760 ;
        RECT 62.860 225.065 62.870 225.760 ;
        RECT 66.540 225.065 66.550 225.760 ;
        RECT 70.220 225.065 70.230 225.760 ;
        RECT 73.900 225.065 73.910 225.760 ;
        RECT 77.580 225.065 77.590 225.760 ;
        RECT 81.260 225.065 81.270 225.760 ;
        RECT 84.940 225.065 84.950 225.760 ;
        RECT 88.620 225.065 88.630 225.760 ;
        RECT 3.480 224.760 3.990 225.065 ;
        RECT 4.290 224.765 7.670 225.065 ;
        RECT 7.970 224.765 11.350 225.065 ;
        RECT 11.650 224.765 15.030 225.065 ;
        RECT 15.330 224.765 18.710 225.065 ;
        RECT 19.010 224.765 22.390 225.065 ;
        RECT 22.690 224.765 26.070 225.065 ;
        RECT 26.370 224.765 29.750 225.065 ;
        RECT 30.050 224.765 33.430 225.065 ;
        RECT 33.730 224.765 37.110 225.065 ;
        RECT 37.410 224.765 40.790 225.065 ;
        RECT 41.090 224.765 44.470 225.065 ;
        RECT 44.770 224.765 48.150 225.065 ;
        RECT 48.450 224.765 51.830 225.065 ;
        RECT 52.130 224.765 55.510 225.065 ;
        RECT 55.810 224.765 59.190 225.065 ;
        RECT 59.490 224.765 62.870 225.065 ;
        RECT 63.170 224.765 66.550 225.065 ;
        RECT 66.850 224.765 70.230 225.065 ;
        RECT 70.530 224.765 73.910 225.065 ;
        RECT 74.210 224.765 77.590 225.065 ;
        RECT 77.890 224.765 81.270 225.065 ;
        RECT 81.570 224.765 84.950 225.065 ;
        RECT 85.250 224.765 88.630 225.065 ;
        RECT 92.300 224.770 92.310 225.760 ;
        RECT 95.980 224.770 95.990 225.760 ;
        RECT 99.660 224.770 99.670 225.760 ;
        RECT 103.340 224.770 103.350 225.760 ;
        RECT 107.020 224.770 107.030 225.760 ;
        RECT 110.700 224.770 110.710 225.760 ;
        RECT 114.380 224.770 114.390 225.760 ;
        RECT 118.060 224.770 118.070 225.760 ;
        RECT 121.740 224.770 121.750 225.760 ;
        RECT 125.420 224.770 125.430 225.760 ;
        RECT 129.100 224.770 129.110 225.760 ;
        RECT 132.780 224.770 132.790 225.760 ;
        RECT 136.460 224.770 136.470 225.760 ;
        RECT 140.140 224.770 140.150 225.760 ;
        RECT 143.820 224.770 143.830 225.760 ;
        RECT 147.500 224.770 147.510 225.760 ;
        RECT 151.180 224.770 151.190 225.760 ;
        RECT 154.860 224.770 154.870 225.760 ;
        RECT 158.540 224.770 158.550 225.760 ;
        RECT 4.290 224.760 5.480 224.765 ;
        RECT 3.480 148.665 5.480 224.760 ;
        RECT 17.635 148.665 19.965 148.810 ;
        RECT 3.480 146.665 20.075 148.665 ;
        RECT 143.725 147.680 146.055 147.825 ;
        RECT 158.345 147.680 160.345 224.160 ;
        RECT 3.480 54.905 5.480 146.665 ;
        RECT 17.635 146.480 19.965 146.665 ;
        RECT 143.725 145.680 160.345 147.680 ;
        RECT 143.725 145.495 146.055 145.680 ;
        RECT 100.595 60.195 101.325 60.925 ;
        RECT 3.480 54.895 4.585 54.905 ;
        RECT 4.595 54.895 5.480 54.905 ;
        RECT 3.480 29.585 5.480 54.895 ;
        RECT 70.945 54.185 72.075 55.315 ;
        RECT 71.360 52.280 71.660 54.185 ;
        RECT 57.560 51.980 71.660 52.280 ;
        RECT 57.560 43.755 57.860 51.980 ;
        RECT 71.360 51.565 71.660 51.980 ;
        RECT 70.945 50.435 72.075 51.565 ;
        RECT 55.940 43.735 57.860 43.755 ;
        RECT 54.925 43.455 57.860 43.735 ;
        RECT 54.925 43.435 56.240 43.455 ;
        RECT 54.925 31.950 55.225 43.435 ;
        RECT 100.610 34.630 101.310 60.195 ;
        RECT 158.345 43.415 160.345 145.680 ;
        RECT 158.345 43.405 159.280 43.415 ;
        RECT 159.290 43.405 160.345 43.415 ;
        RECT 55.880 31.950 56.610 32.165 ;
        RECT 54.925 31.650 56.610 31.950 ;
        RECT 55.880 31.435 56.610 31.650 ;
        RECT 17.635 29.585 19.965 29.730 ;
        RECT 3.480 27.585 20.075 29.585 ;
        RECT 3.480 1.015 5.480 27.585 ;
        RECT 17.635 27.400 19.965 27.585 ;
        RECT 100.230 12.460 122.405 34.630 ;
        RECT 143.725 16.850 146.055 16.995 ;
        RECT 158.345 16.850 160.345 43.405 ;
        RECT 143.725 14.850 160.345 16.850 ;
        RECT 143.725 14.665 146.055 14.850 ;
        RECT 144.890 10.355 157.725 10.590 ;
        RECT 144.125 8.825 157.725 10.355 ;
        RECT 144.890 8.590 157.725 8.825 ;
        RECT 133.795 6.615 135.325 8.145 ;
        RECT 111.860 4.695 113.390 6.225 ;
        RECT 89.520 4.290 91.050 4.560 ;
        RECT 67.345 2.960 68.875 3.055 ;
        RECT 89.520 3.030 91.150 4.290 ;
        RECT 67.345 1.525 69.005 2.960 ;
        RECT 1.990 1.000 2.590 1.010 ;
        RECT 24.070 1.000 24.670 1.010 ;
        RECT 46.150 1.000 46.750 1.010 ;
        RECT 68.005 1.000 69.005 1.525 ;
        RECT 1.990 0.010 2.000 1.000 ;
        RECT 24.070 0.010 24.080 1.000 ;
        RECT 46.150 0.010 46.160 1.000 ;
        RECT 68.005 0.680 68.240 1.000 ;
        RECT 68.840 0.680 69.005 1.000 ;
        RECT 90.150 1.000 91.150 3.030 ;
        RECT 90.150 0.840 90.320 1.000 ;
        RECT 90.920 0.840 91.150 1.000 ;
        RECT 112.130 1.000 113.130 4.695 ;
        RECT 68.230 0.010 68.240 0.680 ;
        RECT 90.310 0.010 90.320 0.840 ;
        RECT 112.130 0.505 112.400 1.000 ;
        RECT 113.000 0.505 113.130 1.000 ;
        RECT 134.280 1.000 135.280 6.615 ;
        RECT 134.280 0.800 134.480 1.000 ;
        RECT 135.080 0.800 135.280 1.000 ;
        RECT 155.725 1.000 157.725 8.590 ;
        RECT 158.345 1.015 160.345 14.850 ;
        RECT 112.390 0.010 112.400 0.505 ;
        RECT 134.470 0.010 134.480 0.800 ;
        RECT 155.725 0.680 156.560 1.000 ;
        RECT 157.160 0.680 157.725 1.000 ;
        RECT 156.550 0.010 156.560 0.680 ;
  END
END tt_um_Burrows_Katie
END LIBRARY

