VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OpAmp
  CLASS BLOCK ;
  FOREIGN OpAmp ;
  ORIGIN 0.000 100.255 ;
  SIZE 99.805 BY 100.255 ;
  PIN VDD
    ANTENNADIFFAREA 133.070694 ;
    PORT
      LAYER nwell ;
        RECT 16.205 -15.170 29.175 -8.750 ;
        RECT 34.740 -15.165 47.710 -8.745 ;
        RECT 54.400 -17.980 66.740 -9.560 ;
        RECT 16.205 -33.515 29.175 -27.095 ;
        RECT 34.495 -33.820 47.465 -27.400 ;
        RECT 2.910 -56.915 8.190 -50.495 ;
        RECT 12.800 -56.915 18.080 -50.495 ;
        RECT 22.635 -56.960 27.915 -50.540 ;
        RECT 32.195 -56.915 37.475 -50.495 ;
        RECT 41.720 -54.645 55.520 -46.225 ;
        RECT 59.365 -54.625 73.165 -46.205 ;
        RECT 2.865 -66.195 8.145 -59.775 ;
        RECT 12.740 -66.195 18.020 -59.775 ;
        RECT 22.680 -66.195 27.960 -59.775 ;
        RECT 32.100 -66.195 37.380 -59.775 ;
        RECT 42.200 -67.000 55.940 -58.580 ;
        RECT 58.905 -66.745 72.645 -58.325 ;
        RECT 2.865 -76.345 8.145 -69.925 ;
        RECT 12.760 -76.345 18.040 -69.925 ;
        RECT 22.805 -76.345 28.085 -69.925 ;
        RECT 32.005 -76.345 37.285 -69.925 ;
      LAYER li1 ;
        RECT 11.310 -7.055 11.980 -6.885 ;
        RECT 21.915 -8.970 22.615 -7.855 ;
        RECT 40.520 -8.965 41.220 -8.130 ;
        RECT 16.540 -9.300 28.840 -8.970 ;
        RECT 35.075 -9.295 47.375 -8.965 ;
        RECT 59.850 -9.780 60.550 -8.405 ;
        RECT 54.735 -10.110 66.405 -9.780 ;
        RECT 54.815 -16.060 54.985 -10.525 ;
        RECT 53.655 -16.760 54.985 -16.060 ;
        RECT 54.815 -17.315 54.985 -16.760 ;
        RECT 56.075 -18.700 56.245 -10.525 ;
        RECT 54.830 -18.870 56.245 -18.700 ;
        RECT 54.830 -19.865 55.000 -18.870 ;
        RECT 57.335 -19.640 57.505 -10.525 ;
        RECT 53.655 -20.035 55.000 -19.865 ;
        RECT 55.865 -19.810 57.505 -19.640 ;
        RECT 53.655 -20.645 53.825 -20.035 ;
        RECT 55.865 -20.855 56.035 -19.810 ;
        RECT 58.595 -20.655 58.765 -10.525 ;
        RECT 55.195 -21.025 56.035 -20.855 ;
        RECT 56.970 -20.825 58.765 -20.655 ;
        RECT 55.195 -21.895 55.365 -21.025 ;
        RECT 54.770 -22.065 55.365 -21.895 ;
        RECT 56.970 -22.030 57.140 -20.825 ;
        RECT 54.770 -22.985 54.940 -22.065 ;
        RECT 53.655 -23.155 54.940 -22.985 ;
        RECT 56.730 -22.200 57.140 -22.030 ;
        RECT 59.855 -22.100 60.025 -10.525 ;
        RECT 56.730 -23.095 56.900 -22.200 ;
        RECT 58.900 -22.270 60.025 -22.100 ;
        RECT 61.115 -22.260 61.285 -10.525 ;
        RECT 62.375 -20.760 62.545 -10.525 ;
        RECT 63.635 -19.650 63.805 -10.525 ;
        RECT 64.895 -18.600 65.065 -10.525 ;
        RECT 66.155 -16.325 66.325 -10.525 ;
        RECT 67.125 -16.325 67.295 -16.145 ;
        RECT 66.155 -16.495 67.295 -16.325 ;
        RECT 66.155 -16.505 66.330 -16.495 ;
        RECT 66.155 -17.315 66.325 -16.505 ;
        RECT 67.125 -16.675 67.295 -16.495 ;
        RECT 64.895 -18.770 66.340 -18.600 ;
        RECT 66.170 -19.445 66.340 -18.770 ;
        RECT 66.170 -19.615 67.525 -19.445 ;
        RECT 63.635 -19.820 65.090 -19.650 ;
        RECT 64.920 -20.475 65.090 -19.820 ;
        RECT 67.355 -19.665 67.525 -19.615 ;
        RECT 67.355 -20.015 67.550 -19.665 ;
        RECT 67.380 -20.195 67.550 -20.015 ;
        RECT 64.920 -20.645 66.090 -20.475 ;
        RECT 62.375 -20.930 63.890 -20.760 ;
        RECT 63.720 -21.555 63.890 -20.930 ;
        RECT 65.920 -21.340 66.090 -20.645 ;
        RECT 65.920 -21.510 66.525 -21.340 ;
        RECT 63.720 -21.725 64.395 -21.555 ;
        RECT 53.655 -23.650 53.825 -23.155 ;
        RECT 58.900 -23.605 59.070 -22.270 ;
        RECT 61.115 -22.430 62.350 -22.260 ;
        RECT 62.180 -23.605 62.350 -22.430 ;
        RECT 64.225 -23.095 64.395 -21.725 ;
        RECT 66.355 -22.430 66.525 -21.510 ;
        RECT 66.355 -22.600 67.535 -22.430 ;
        RECT 67.355 -22.915 67.535 -22.600 ;
        RECT 67.355 -23.095 67.525 -22.915 ;
        RECT 58.900 -23.955 59.075 -23.605 ;
        RECT 62.180 -23.955 62.355 -23.605 ;
        RECT 58.905 -24.135 59.075 -23.955 ;
        RECT 62.185 -24.135 62.355 -23.955 ;
        RECT 17.345 -26.265 18.345 -25.265 ;
        RECT 17.785 -27.315 18.115 -26.265 ;
        RECT 45.960 -26.760 46.490 -26.230 ;
        RECT 16.540 -27.645 28.840 -27.315 ;
        RECT 46.075 -27.620 46.375 -26.760 ;
        RECT 34.830 -27.950 47.130 -27.620 ;
        RECT 57.415 -46.440 57.945 -46.335 ;
        RECT 59.700 -46.440 72.830 -46.425 ;
        RECT 42.055 -46.470 55.185 -46.445 ;
        RECT 57.245 -46.470 72.830 -46.440 ;
        RECT 42.055 -46.755 72.830 -46.470 ;
        RECT 42.055 -46.770 59.910 -46.755 ;
        RECT 42.055 -46.775 55.185 -46.770 ;
        RECT 57.415 -46.865 57.945 -46.770 ;
        RECT 3.245 -51.045 9.145 -50.715 ;
        RECT 13.135 -51.045 18.660 -50.715 ;
        RECT 8.815 -51.330 9.145 -51.045 ;
        RECT 18.330 -51.330 18.660 -51.045 ;
        RECT 22.970 -50.935 28.900 -50.760 ;
        RECT 22.970 -51.090 28.905 -50.935 ;
        RECT 32.530 -51.045 38.505 -50.715 ;
        RECT 8.860 -51.430 9.030 -51.330 ;
        RECT 18.380 -51.430 18.550 -51.330 ;
        RECT 28.735 -51.465 28.905 -51.090 ;
        RECT 38.175 -51.335 38.505 -51.045 ;
        RECT 31.905 -51.475 32.075 -51.465 ;
        RECT 3.325 -51.495 3.495 -51.480 ;
        RECT 13.215 -51.495 13.385 -51.480 ;
        RECT 1.895 -52.195 3.505 -51.495 ;
        RECT 11.800 -52.195 13.410 -51.495 ;
        RECT 23.050 -51.545 23.220 -51.525 ;
        RECT 3.325 -56.230 3.495 -52.195 ;
        RECT 13.215 -56.230 13.385 -52.195 ;
        RECT 21.610 -52.245 23.220 -51.545 ;
        RECT 31.905 -51.995 32.795 -51.475 ;
        RECT 31.910 -52.175 32.795 -51.995 ;
        RECT 23.050 -56.275 23.220 -52.245 ;
        RECT 32.610 -56.230 32.780 -52.175 ;
        RECT 42.135 -54.670 42.305 -47.190 ;
        RECT 44.695 -54.670 44.865 -47.190 ;
        RECT 47.255 -54.670 47.425 -47.190 ;
        RECT 49.815 -54.670 49.985 -47.190 ;
        RECT 52.375 -54.670 52.545 -47.190 ;
        RECT 54.935 -54.670 55.105 -47.190 ;
        RECT 59.780 -53.780 59.950 -47.170 ;
        RECT 59.780 -53.960 59.955 -53.780 ;
        RECT 62.340 -53.890 62.510 -47.170 ;
        RECT 64.900 -53.890 65.070 -47.170 ;
        RECT 67.460 -53.890 67.630 -47.170 ;
        RECT 70.020 -53.890 70.190 -47.170 ;
        RECT 72.580 -53.030 72.750 -47.170 ;
        RECT 72.580 -53.200 73.625 -53.030 ;
        RECT 62.340 -53.960 62.515 -53.890 ;
        RECT 64.900 -53.960 65.075 -53.890 ;
        RECT 67.460 -53.960 67.635 -53.890 ;
        RECT 70.020 -53.960 70.195 -53.890 ;
        RECT 72.580 -53.960 72.750 -53.200 ;
        RECT 59.785 -54.670 59.955 -53.960 ;
        RECT 41.960 -55.200 42.490 -54.670 ;
        RECT 44.475 -55.200 45.005 -54.670 ;
        RECT 47.080 -55.200 47.610 -54.670 ;
        RECT 49.610 -55.200 50.140 -54.670 ;
        RECT 52.255 -55.200 52.785 -54.670 ;
        RECT 54.730 -55.200 55.260 -54.670 ;
        RECT 59.605 -55.200 60.135 -54.670 ;
        RECT 62.345 -54.745 62.515 -53.960 ;
        RECT 62.170 -55.275 62.700 -54.745 ;
        RECT 64.905 -54.750 65.075 -53.960 ;
        RECT 67.465 -54.710 67.635 -53.960 ;
        RECT 64.725 -55.280 65.255 -54.750 ;
        RECT 67.290 -55.240 67.820 -54.710 ;
        RECT 70.025 -54.735 70.195 -53.960 ;
        RECT 73.455 -54.260 73.625 -53.200 ;
        RECT 69.850 -55.265 70.380 -54.735 ;
        RECT 73.275 -54.790 73.805 -54.260 ;
        RECT 57.415 -58.545 57.945 -58.490 ;
        RECT 57.415 -58.605 72.310 -58.545 ;
        RECT 5.145 -58.890 5.315 -58.790 ;
        RECT 15.495 -58.890 15.665 -58.790 ;
        RECT 25.355 -58.890 25.525 -58.790 ;
        RECT 5.035 -59.995 5.365 -58.890 ;
        RECT 15.360 -59.995 15.690 -58.890 ;
        RECT 25.300 -59.995 25.630 -58.890 ;
        RECT 34.680 -59.115 34.850 -58.790 ;
        RECT 42.535 -58.850 55.605 -58.800 ;
        RECT 55.870 -58.850 72.310 -58.605 ;
        RECT 42.535 -58.875 72.310 -58.850 ;
        RECT 42.535 -58.905 57.945 -58.875 ;
        RECT 34.630 -59.995 34.960 -59.115 ;
        RECT 42.535 -59.130 56.170 -58.905 ;
        RECT 57.415 -59.020 57.945 -58.905 ;
        RECT 55.370 -59.150 56.170 -59.130 ;
        RECT 3.200 -60.325 7.810 -59.995 ;
        RECT 13.075 -60.325 17.685 -59.995 ;
        RECT 23.015 -60.325 27.625 -59.995 ;
        RECT 32.435 -60.325 37.045 -59.995 ;
        RECT 42.615 -66.215 42.785 -59.545 ;
        RECT 44.435 -66.085 44.605 -59.545 ;
        RECT 42.600 -66.335 42.785 -66.215 ;
        RECT 44.420 -66.335 44.605 -66.085 ;
        RECT 46.255 -66.105 46.425 -59.545 ;
        RECT 46.240 -66.335 46.425 -66.105 ;
        RECT 48.075 -66.215 48.245 -59.545 ;
        RECT 48.060 -66.335 48.245 -66.215 ;
        RECT 42.600 -66.595 42.770 -66.335 ;
        RECT 44.420 -66.595 44.590 -66.335 ;
        RECT 46.240 -66.595 46.410 -66.335 ;
        RECT 42.600 -66.945 42.775 -66.595 ;
        RECT 44.420 -66.945 44.595 -66.595 ;
        RECT 46.240 -66.945 46.415 -66.595 ;
        RECT 42.605 -67.125 42.775 -66.945 ;
        RECT 44.425 -67.125 44.595 -66.945 ;
        RECT 46.245 -67.125 46.415 -66.945 ;
        RECT 48.060 -67.115 48.230 -66.335 ;
        RECT 49.895 -66.585 50.065 -59.545 ;
        RECT 51.715 -66.070 51.885 -59.545 ;
        RECT 49.885 -66.935 50.065 -66.585 ;
        RECT 51.700 -66.335 51.885 -66.070 ;
        RECT 53.535 -66.080 53.705 -59.545 ;
        RECT 53.520 -66.335 53.705 -66.080 ;
        RECT 55.355 -66.120 55.525 -59.545 ;
        RECT 55.340 -66.335 55.525 -66.120 ;
        RECT 51.700 -66.585 51.870 -66.335 ;
        RECT 51.700 -66.935 51.880 -66.585 ;
        RECT 49.885 -67.115 50.055 -66.935 ;
        RECT 51.710 -67.115 51.880 -66.935 ;
        RECT 53.520 -67.125 53.690 -66.335 ;
        RECT 55.340 -66.585 55.510 -66.335 ;
        RECT 55.340 -66.655 55.515 -66.585 ;
        RECT 55.225 -66.850 55.515 -66.655 ;
        RECT 55.345 -67.115 55.515 -66.850 ;
        RECT 5.145 -69.100 5.315 -68.815 ;
        RECT 15.495 -69.055 15.665 -68.815 ;
        RECT 25.515 -69.010 25.685 -68.815 ;
        RECT 5.075 -70.145 5.405 -69.100 ;
        RECT 15.465 -70.145 15.795 -69.055 ;
        RECT 25.450 -70.145 25.780 -69.010 ;
        RECT 34.450 -69.045 34.620 -68.815 ;
        RECT 34.400 -70.145 34.730 -69.045 ;
        RECT 3.200 -70.475 7.810 -70.145 ;
        RECT 13.095 -70.475 17.705 -70.145 ;
        RECT 23.140 -70.475 27.750 -70.145 ;
        RECT 32.340 -70.475 36.950 -70.145 ;
      LAYER met1 ;
        RECT 0.000 -4.880 99.790 0.000 ;
        RECT 3.830 -48.500 4.530 -4.880 ;
        RECT 11.315 -6.960 12.015 -4.880 ;
        RECT 11.320 -7.085 11.970 -6.960 ;
        RECT 12.515 -8.840 13.215 -4.880 ;
        RECT 21.915 -8.975 22.615 -4.880 ;
        RECT 40.520 -8.690 41.220 -4.880 ;
        RECT 17.345 -26.265 18.345 -25.265 ;
        RECT 50.365 -26.115 51.065 -4.880 ;
        RECT 59.810 -9.050 60.510 -4.880 ;
        RECT 66.910 -5.155 67.610 -4.880 ;
        RECT 66.960 -5.520 67.600 -5.155 ;
        RECT 53.420 -15.960 54.060 -15.940 ;
        RECT 66.890 -15.960 67.530 -15.940 ;
        RECT 53.260 -16.860 54.220 -15.960 ;
        RECT 66.730 -16.860 67.690 -15.960 ;
        RECT 53.420 -16.880 54.060 -16.860 ;
        RECT 66.890 -16.880 67.530 -16.860 ;
        RECT 67.145 -19.480 67.785 -19.460 ;
        RECT 53.420 -19.930 54.060 -19.910 ;
        RECT 53.260 -20.830 54.220 -19.930 ;
        RECT 66.985 -20.380 67.945 -19.480 ;
        RECT 67.145 -20.400 67.785 -20.380 ;
        RECT 53.420 -20.850 54.060 -20.830 ;
        RECT 56.495 -22.380 57.135 -22.360 ;
        RECT 63.990 -22.380 64.630 -22.360 ;
        RECT 67.120 -22.380 67.760 -22.360 ;
        RECT 53.420 -22.935 54.060 -22.915 ;
        RECT 53.260 -23.835 54.220 -22.935 ;
        RECT 56.335 -23.280 57.295 -22.380 ;
        RECT 63.830 -23.280 64.790 -22.380 ;
        RECT 66.960 -23.280 67.920 -22.380 ;
        RECT 56.495 -23.300 57.135 -23.280 ;
        RECT 63.990 -23.300 64.630 -23.280 ;
        RECT 67.120 -23.300 67.760 -23.280 ;
        RECT 58.670 -23.420 59.310 -23.400 ;
        RECT 61.950 -23.420 62.590 -23.400 ;
        RECT 53.420 -23.855 54.060 -23.835 ;
        RECT 58.510 -24.320 59.470 -23.420 ;
        RECT 61.790 -24.320 62.750 -23.420 ;
        RECT 58.670 -24.340 59.310 -24.320 ;
        RECT 61.950 -24.340 62.590 -24.320 ;
        RECT 50.365 -26.145 52.435 -26.115 ;
        RECT 46.275 -26.200 52.435 -26.145 ;
        RECT 45.900 -26.790 52.435 -26.200 ;
        RECT 46.275 -26.815 52.435 -26.790 ;
        RECT 46.275 -26.845 51.065 -26.815 ;
        RECT 51.735 -28.600 52.435 -26.815 ;
        RECT 51.735 -29.300 58.030 -28.600 ;
        RECT 3.645 -49.080 4.530 -48.500 ;
        RECT 3.830 -49.125 4.530 -49.080 ;
        RECT 38.020 -50.620 38.660 -50.600 ;
        RECT 8.625 -50.715 9.265 -50.695 ;
        RECT 18.145 -50.715 18.785 -50.695 ;
        RECT 1.715 -51.365 2.355 -51.345 ;
        RECT 1.555 -52.265 2.515 -51.365 ;
        RECT 8.465 -51.615 9.425 -50.715 ;
        RECT 11.715 -51.440 12.355 -51.420 ;
        RECT 8.625 -51.635 9.265 -51.615 ;
        RECT 1.715 -52.285 2.355 -52.265 ;
        RECT 11.555 -52.340 12.515 -51.440 ;
        RECT 17.985 -51.615 18.945 -50.715 ;
        RECT 28.500 -50.750 29.140 -50.730 ;
        RECT 21.545 -51.440 22.185 -51.420 ;
        RECT 18.145 -51.635 18.785 -51.615 ;
        RECT 21.385 -52.340 22.345 -51.440 ;
        RECT 28.340 -51.650 29.300 -50.750 ;
        RECT 31.670 -51.280 32.310 -51.260 ;
        RECT 28.500 -51.670 29.140 -51.650 ;
        RECT 31.510 -52.180 32.470 -51.280 ;
        RECT 37.860 -51.520 38.820 -50.620 ;
        RECT 38.020 -51.540 38.660 -51.520 ;
        RECT 31.670 -52.200 32.310 -52.180 ;
        RECT 11.715 -52.360 12.355 -52.340 ;
        RECT 21.545 -52.360 22.185 -52.340 ;
        RECT 57.330 -54.585 58.030 -29.300 ;
        RECT 59.800 -54.585 59.940 -54.470 ;
        RECT 41.900 -54.865 42.550 -54.640 ;
        RECT 44.415 -54.865 45.065 -54.640 ;
        RECT 47.020 -54.865 47.670 -54.640 ;
        RECT 49.550 -54.865 50.200 -54.640 ;
        RECT 52.195 -54.865 52.845 -54.640 ;
        RECT 54.670 -54.865 55.320 -54.640 ;
        RECT 41.900 -55.005 55.320 -54.865 ;
        RECT 41.900 -55.230 42.550 -55.005 ;
        RECT 44.415 -55.230 45.065 -55.005 ;
        RECT 47.020 -55.230 47.670 -55.005 ;
        RECT 49.550 -55.230 50.200 -55.005 ;
        RECT 52.195 -55.230 52.845 -55.005 ;
        RECT 54.670 -55.230 55.320 -55.005 ;
        RECT 57.330 -54.940 60.220 -54.585 ;
        RECT 62.110 -54.940 62.760 -54.715 ;
        RECT 57.330 -54.945 62.760 -54.940 ;
        RECT 64.665 -54.905 65.315 -54.720 ;
        RECT 67.230 -54.905 67.880 -54.680 ;
        RECT 64.665 -54.930 67.880 -54.905 ;
        RECT 69.790 -54.930 70.440 -54.705 ;
        RECT 73.215 -54.820 73.865 -54.230 ;
        RECT 64.665 -54.945 70.440 -54.930 ;
        RECT 57.330 -54.985 70.440 -54.945 ;
        RECT 73.470 -54.985 73.610 -54.820 ;
        RECT 57.330 -55.045 73.610 -54.985 ;
        RECT 57.330 -55.080 65.315 -55.045 ;
        RECT 42.155 -55.910 42.295 -55.230 ;
        RECT 57.330 -55.285 60.220 -55.080 ;
        RECT 41.905 -56.490 42.545 -55.910 ;
        RECT 4.910 -58.605 5.550 -58.585 ;
        RECT 15.260 -58.605 15.900 -58.585 ;
        RECT 25.120 -58.605 25.760 -58.585 ;
        RECT 34.445 -58.605 35.085 -58.585 ;
        RECT 4.750 -59.505 5.710 -58.605 ;
        RECT 15.100 -59.505 16.060 -58.605 ;
        RECT 24.960 -59.505 25.920 -58.605 ;
        RECT 34.285 -59.505 35.245 -58.605 ;
        RECT 57.330 -59.050 58.030 -55.285 ;
        RECT 59.520 -55.345 60.220 -55.285 ;
        RECT 62.110 -55.085 65.315 -55.080 ;
        RECT 62.110 -55.305 62.760 -55.085 ;
        RECT 64.665 -55.310 65.315 -55.085 ;
        RECT 67.230 -55.070 73.610 -55.045 ;
        RECT 67.230 -55.270 67.880 -55.070 ;
        RECT 69.790 -55.125 73.610 -55.070 ;
        RECT 69.790 -55.295 70.440 -55.125 ;
        RECT 4.910 -59.525 5.550 -59.505 ;
        RECT 15.260 -59.525 15.900 -59.505 ;
        RECT 25.120 -59.525 25.760 -59.505 ;
        RECT 34.445 -59.525 35.085 -59.505 ;
        RECT 42.370 -66.410 43.010 -66.390 ;
        RECT 44.190 -66.410 44.830 -66.390 ;
        RECT 46.010 -66.410 46.650 -66.390 ;
        RECT 47.825 -66.400 48.465 -66.380 ;
        RECT 49.650 -66.400 50.290 -66.380 ;
        RECT 51.475 -66.400 52.115 -66.380 ;
        RECT 42.210 -67.310 43.170 -66.410 ;
        RECT 44.030 -67.310 44.990 -66.410 ;
        RECT 45.850 -67.310 46.810 -66.410 ;
        RECT 47.665 -67.300 48.625 -66.400 ;
        RECT 49.490 -67.300 50.450 -66.400 ;
        RECT 51.315 -67.300 52.275 -66.400 ;
        RECT 53.285 -66.410 53.925 -66.390 ;
        RECT 55.110 -66.400 55.750 -66.380 ;
        RECT 42.370 -67.330 43.010 -67.310 ;
        RECT 44.190 -67.330 44.830 -67.310 ;
        RECT 46.010 -67.330 46.650 -67.310 ;
        RECT 47.825 -67.320 48.465 -67.300 ;
        RECT 49.650 -67.320 50.290 -67.300 ;
        RECT 51.475 -67.320 52.115 -67.300 ;
        RECT 53.125 -67.310 54.085 -66.410 ;
        RECT 54.950 -67.300 55.910 -66.400 ;
        RECT 53.285 -67.330 53.925 -67.310 ;
        RECT 55.110 -67.320 55.750 -67.300 ;
        RECT 4.910 -68.630 5.550 -68.610 ;
        RECT 15.260 -68.630 15.900 -68.610 ;
        RECT 25.280 -68.630 25.920 -68.610 ;
        RECT 34.215 -68.630 34.855 -68.610 ;
        RECT 4.750 -69.530 5.710 -68.630 ;
        RECT 15.100 -69.530 16.060 -68.630 ;
        RECT 25.120 -69.530 26.080 -68.630 ;
        RECT 34.055 -69.530 35.015 -68.630 ;
        RECT 4.910 -69.550 5.550 -69.530 ;
        RECT 15.260 -69.550 15.900 -69.530 ;
        RECT 25.280 -69.550 25.920 -69.530 ;
        RECT 34.215 -69.550 34.855 -69.530 ;
      LAYER met2 ;
        RECT 66.960 -5.155 67.600 -4.930 ;
        RECT 12.480 -8.905 13.250 -8.175 ;
        RECT 66.910 -15.960 67.610 -5.155 ;
        RECT 53.260 -16.060 54.220 -15.960 ;
        RECT 52.030 -16.760 54.220 -16.060 ;
        RECT 52.030 -20.005 52.730 -16.760 ;
        RECT 53.260 -16.860 54.220 -16.760 ;
        RECT 66.730 -16.060 67.690 -15.960 ;
        RECT 66.730 -16.760 69.395 -16.060 ;
        RECT 66.730 -16.860 67.690 -16.760 ;
        RECT 66.985 -19.615 67.945 -19.480 ;
        RECT 68.695 -19.615 69.395 -16.760 ;
        RECT 53.260 -20.005 54.220 -19.930 ;
        RECT 52.030 -20.705 54.220 -20.005 ;
        RECT 66.985 -20.315 69.395 -19.615 ;
        RECT 66.985 -20.380 67.945 -20.315 ;
        RECT 52.030 -23.035 52.730 -20.705 ;
        RECT 53.260 -20.830 54.220 -20.705 ;
        RECT 53.260 -23.035 54.220 -22.935 ;
        RECT 52.030 -23.735 54.220 -23.035 ;
        RECT 56.335 -23.080 59.015 -22.380 ;
        RECT 56.335 -23.280 57.295 -23.080 ;
        RECT 53.260 -23.835 54.220 -23.735 ;
        RECT 58.315 -23.420 59.015 -23.080 ;
        RECT 63.830 -22.760 64.790 -22.380 ;
        RECT 66.960 -22.760 67.920 -22.380 ;
        RECT 68.695 -22.425 69.395 -20.315 ;
        RECT 63.830 -22.775 67.920 -22.760 ;
        RECT 68.450 -22.775 69.395 -22.425 ;
        RECT 63.830 -22.845 69.395 -22.775 ;
        RECT 63.830 -22.900 69.150 -22.845 ;
        RECT 63.830 -23.280 64.790 -22.900 ;
        RECT 66.960 -22.915 69.150 -22.900 ;
        RECT 66.960 -23.280 67.920 -22.915 ;
        RECT 17.260 -26.330 18.430 -25.200 ;
        RECT 53.390 -25.565 54.090 -23.835 ;
        RECT 58.315 -24.220 59.470 -23.420 ;
        RECT 58.510 -24.320 59.470 -24.220 ;
        RECT 61.790 -24.320 62.750 -23.420 ;
        RECT 58.640 -25.565 59.340 -24.320 ;
        RECT 53.390 -25.625 59.340 -25.565 ;
        RECT 61.920 -25.625 62.620 -24.320 ;
        RECT 53.390 -25.640 62.825 -25.625 ;
        RECT 68.450 -25.640 69.150 -22.915 ;
        RECT 53.390 -26.265 69.150 -25.640 ;
        RECT 58.640 -26.325 69.150 -26.265 ;
        RECT 62.125 -26.340 69.150 -26.325 ;
        RECT 3.570 -49.140 4.285 -48.440 ;
        RECT 3.570 -49.310 4.270 -49.140 ;
        RECT 1.615 -50.010 40.950 -49.310 ;
        RECT 1.615 -51.365 2.315 -50.010 ;
        RECT 8.465 -50.930 9.425 -50.715 ;
        RECT 9.565 -50.930 10.265 -50.010 ;
        RECT 1.555 -52.265 2.515 -51.365 ;
        RECT 8.465 -51.570 10.265 -50.930 ;
        RECT 17.985 -50.815 18.945 -50.715 ;
        RECT 19.840 -50.815 20.540 -50.010 ;
        RECT 11.555 -51.570 12.515 -51.440 ;
        RECT 8.465 -51.615 12.515 -51.570 ;
        RECT 17.985 -51.515 20.540 -50.815 ;
        RECT 28.340 -50.775 29.300 -50.750 ;
        RECT 30.035 -50.775 30.735 -50.010 ;
        RECT 28.340 -51.410 30.735 -50.775 ;
        RECT 37.860 -50.655 38.820 -50.620 ;
        RECT 40.250 -50.655 40.950 -50.010 ;
        RECT 31.510 -51.410 32.470 -51.280 ;
        RECT 17.985 -51.615 18.945 -51.515 ;
        RECT 19.840 -51.595 20.540 -51.515 ;
        RECT 21.385 -51.595 22.345 -51.440 ;
        RECT 8.595 -51.630 12.515 -51.615 ;
        RECT 9.565 -52.270 12.515 -51.630 ;
        RECT 11.555 -52.340 12.515 -52.270 ;
        RECT 19.840 -52.295 22.345 -51.595 ;
        RECT 28.340 -51.475 32.470 -51.410 ;
        RECT 28.340 -51.650 29.300 -51.475 ;
        RECT 30.035 -52.110 32.470 -51.475 ;
        RECT 37.860 -51.355 40.950 -50.655 ;
        RECT 37.860 -51.520 38.820 -51.355 ;
        RECT 31.510 -52.180 32.470 -52.110 ;
        RECT 21.385 -52.340 22.345 -52.295 ;
        RECT 40.250 -55.850 40.950 -51.355 ;
        RECT 40.250 -56.550 42.545 -55.850 ;
        RECT 4.750 -58.705 5.710 -58.605 ;
        RECT 15.100 -58.705 16.060 -58.605 ;
        RECT 24.960 -58.705 25.920 -58.605 ;
        RECT 34.285 -58.705 35.245 -58.605 ;
        RECT 40.250 -58.705 40.950 -56.550 ;
        RECT 4.750 -59.405 40.950 -58.705 ;
        RECT 4.750 -59.505 5.710 -59.405 ;
        RECT 15.100 -59.505 16.060 -59.405 ;
        RECT 24.960 -59.505 25.920 -59.405 ;
        RECT 34.285 -59.505 35.245 -59.405 ;
        RECT 40.250 -67.785 40.950 -59.405 ;
        RECT 42.210 -67.310 43.170 -66.410 ;
        RECT 44.030 -67.310 44.990 -66.410 ;
        RECT 45.850 -67.310 46.810 -66.410 ;
        RECT 47.665 -67.300 48.625 -66.400 ;
        RECT 49.490 -67.300 50.450 -66.400 ;
        RECT 51.315 -67.300 52.275 -66.400 ;
        RECT 42.620 -67.785 42.760 -67.310 ;
        RECT 44.590 -67.785 44.730 -67.310 ;
        RECT 46.240 -67.785 46.380 -67.310 ;
        RECT 48.105 -67.785 48.245 -67.300 ;
        RECT 49.910 -67.785 50.050 -67.300 ;
        RECT 51.735 -67.785 51.875 -67.300 ;
        RECT 53.125 -67.310 54.085 -66.410 ;
        RECT 54.950 -67.300 55.910 -66.400 ;
        RECT 53.660 -67.785 53.800 -67.310 ;
        RECT 55.285 -67.785 55.425 -67.300 ;
        RECT 40.250 -67.925 55.425 -67.785 ;
        RECT 4.750 -68.850 5.710 -68.630 ;
        RECT 15.100 -68.850 16.060 -68.630 ;
        RECT 25.120 -68.850 26.080 -68.630 ;
        RECT 34.055 -68.850 35.015 -68.630 ;
        RECT 40.250 -68.850 40.950 -67.925 ;
        RECT 4.750 -69.530 40.950 -68.850 ;
        RECT 4.880 -69.550 40.950 -69.530 ;
      LAYER met3 ;
        RECT 12.480 -8.905 13.250 -8.175 ;
        RECT 12.515 -25.455 13.215 -8.905 ;
        RECT 17.260 -25.455 18.430 -25.200 ;
        RECT 12.515 -26.155 18.430 -25.455 ;
        RECT 17.260 -26.330 18.430 -26.155 ;
    END
  END VDD
  PIN Vss
    ANTENNADIFFAREA 51.520798 ;
    PORT
      LAYER pwell ;
        RECT 76.095 -58.245 77.515 -50.975 ;
        RECT 76.015 -58.915 77.595 -58.245 ;
        RECT 76.270 -71.695 77.690 -64.425 ;
        RECT 76.190 -72.365 77.770 -71.695 ;
        RECT 40.420 -79.255 44.210 -72.985 ;
        RECT 47.110 -79.255 50.900 -72.985 ;
        RECT 53.800 -79.255 57.590 -72.985 ;
        RECT 60.440 -79.255 64.230 -72.985 ;
        RECT 3.165 -84.940 7.955 -79.670 ;
        RECT 12.980 -84.940 17.770 -79.670 ;
        RECT 23.140 -84.940 27.930 -79.670 ;
        RECT 32.205 -84.940 36.995 -79.670 ;
        RECT 40.340 -79.925 44.290 -79.255 ;
        RECT 47.030 -79.925 50.980 -79.255 ;
        RECT 53.720 -79.925 57.670 -79.255 ;
        RECT 60.360 -79.925 64.310 -79.255 ;
        RECT 66.640 -82.600 70.430 -76.230 ;
        RECT 73.335 -82.600 77.125 -76.230 ;
        RECT 79.450 -82.600 83.240 -76.230 ;
        RECT 85.855 -82.600 89.645 -76.230 ;
        RECT 66.560 -83.270 70.510 -82.600 ;
        RECT 73.255 -83.270 77.205 -82.600 ;
        RECT 79.370 -83.270 83.320 -82.600 ;
        RECT 85.775 -83.270 89.725 -82.600 ;
        RECT 3.085 -85.610 8.035 -84.940 ;
        RECT 12.900 -85.610 17.850 -84.940 ;
        RECT 23.060 -85.610 28.010 -84.940 ;
        RECT 32.125 -85.610 37.075 -84.940 ;
        RECT 66.640 -92.725 70.430 -86.355 ;
        RECT 73.335 -92.725 77.125 -86.355 ;
        RECT 79.450 -92.725 83.240 -86.355 ;
        RECT 85.855 -92.725 89.645 -86.355 ;
        RECT 66.560 -93.395 70.510 -92.725 ;
        RECT 73.255 -93.395 77.205 -92.725 ;
        RECT 79.370 -93.395 83.320 -92.725 ;
        RECT 85.775 -93.395 89.725 -92.725 ;
      LAYER li1 ;
        RECT 76.185 -58.745 77.425 -58.415 ;
        RECT 76.655 -59.815 76.985 -58.745 ;
        RECT 76.715 -59.915 76.885 -59.815 ;
        RECT 83.315 -67.335 83.985 -67.165 ;
        RECT 76.360 -72.195 77.600 -71.865 ;
        RECT 76.405 -72.465 76.735 -72.195 ;
        RECT 74.720 -72.795 76.735 -72.465 ;
        RECT 74.720 -72.995 75.050 -72.795 ;
        RECT 39.635 -78.690 39.805 -78.590 ;
        RECT 39.540 -78.820 39.870 -78.690 ;
        RECT 40.590 -78.820 40.760 -73.230 ;
        RECT 46.175 -78.690 46.345 -78.590 ;
        RECT 39.540 -78.990 40.760 -78.820 ;
        RECT 39.540 -79.425 39.870 -78.990 ;
        RECT 40.590 -79.000 40.760 -78.990 ;
        RECT 46.145 -78.830 46.475 -78.690 ;
        RECT 47.280 -78.830 47.450 -73.230 ;
        RECT 52.870 -78.690 53.040 -78.590 ;
        RECT 46.145 -79.000 47.450 -78.830 ;
        RECT 52.800 -78.825 53.130 -78.690 ;
        RECT 53.970 -78.825 54.140 -73.230 ;
        RECT 52.800 -78.995 54.140 -78.825 ;
        RECT 46.145 -79.425 46.475 -79.000 ;
        RECT 52.800 -79.425 53.130 -78.995 ;
        RECT 53.970 -79.000 54.140 -78.995 ;
        RECT 59.600 -78.830 59.970 -78.665 ;
        RECT 60.610 -78.830 60.780 -73.230 ;
        RECT 59.600 -79.000 60.780 -78.830 ;
        RECT 59.600 -79.195 59.970 -79.000 ;
        RECT 59.600 -79.425 59.930 -79.195 ;
        RECT 39.540 -79.755 44.120 -79.425 ;
        RECT 46.145 -79.755 50.810 -79.425 ;
        RECT 52.800 -79.755 57.500 -79.425 ;
        RECT 59.600 -79.755 64.140 -79.425 ;
        RECT 2.485 -84.460 2.655 -84.275 ;
        RECT 3.335 -84.460 3.505 -79.925 ;
        RECT 11.335 -84.460 11.505 -84.275 ;
        RECT 13.150 -84.460 13.320 -79.925 ;
        RECT 2.485 -84.630 3.510 -84.460 ;
        RECT 11.335 -84.630 13.320 -84.460 ;
        RECT 2.485 -84.805 2.655 -84.630 ;
        RECT 3.335 -84.675 3.505 -84.630 ;
        RECT 11.335 -84.805 11.505 -84.630 ;
        RECT 13.150 -84.675 13.320 -84.630 ;
        RECT 22.555 -84.460 22.725 -84.275 ;
        RECT 23.310 -84.460 23.480 -79.925 ;
        RECT 22.555 -84.630 23.480 -84.460 ;
        RECT 22.555 -84.805 22.725 -84.630 ;
        RECT 23.310 -84.675 23.480 -84.630 ;
        RECT 31.630 -84.460 31.800 -84.275 ;
        RECT 32.375 -84.460 32.545 -79.925 ;
        RECT 66.105 -82.110 66.275 -81.925 ;
        RECT 66.810 -82.110 66.980 -76.525 ;
        RECT 72.735 -82.110 72.905 -81.925 ;
        RECT 73.505 -82.110 73.675 -76.525 ;
        RECT 78.895 -80.920 79.065 -80.735 ;
        RECT 79.620 -80.920 79.790 -76.525 ;
        RECT 78.895 -81.090 79.790 -80.920 ;
        RECT 78.895 -81.265 79.065 -81.090 ;
        RECT 66.105 -82.280 66.995 -82.110 ;
        RECT 72.735 -82.280 73.675 -82.110 ;
        RECT 66.105 -82.455 66.275 -82.280 ;
        RECT 66.810 -82.295 66.980 -82.280 ;
        RECT 72.735 -82.455 72.905 -82.280 ;
        RECT 73.505 -82.295 73.675 -82.280 ;
        RECT 79.620 -82.295 79.790 -81.090 ;
        RECT 85.300 -80.920 85.470 -80.735 ;
        RECT 86.025 -80.920 86.195 -76.525 ;
        RECT 85.300 -81.090 86.195 -80.920 ;
        RECT 85.300 -81.265 85.470 -81.090 ;
        RECT 86.025 -82.295 86.195 -81.090 ;
        RECT 66.730 -83.100 70.340 -82.770 ;
        RECT 73.425 -83.100 77.035 -82.770 ;
        RECT 79.540 -83.100 83.150 -82.770 ;
        RECT 85.945 -83.100 89.555 -82.770 ;
        RECT 68.130 -83.855 68.460 -83.100 ;
        RECT 75.175 -83.855 75.505 -83.100 ;
        RECT 68.245 -83.955 68.415 -83.855 ;
        RECT 75.210 -83.955 75.380 -83.855 ;
        RECT 81.415 -83.955 81.745 -83.100 ;
        RECT 87.500 -83.855 87.830 -83.100 ;
        RECT 87.570 -83.955 87.740 -83.855 ;
        RECT 31.630 -84.630 32.545 -84.460 ;
        RECT 31.630 -84.805 31.800 -84.630 ;
        RECT 32.375 -84.675 32.545 -84.630 ;
        RECT 3.255 -85.440 7.865 -85.110 ;
        RECT 13.070 -85.440 17.680 -85.110 ;
        RECT 23.230 -85.440 27.840 -85.110 ;
        RECT 32.295 -85.440 36.905 -85.110 ;
        RECT 4.500 -86.795 5.500 -85.440 ;
        RECT 14.295 -86.795 15.295 -85.440 ;
        RECT 23.655 -86.795 24.655 -85.440 ;
        RECT 34.225 -87.165 35.225 -85.440 ;
        RECT 66.100 -86.685 66.270 -86.500 ;
        RECT 66.810 -86.685 66.980 -86.650 ;
        RECT 72.760 -86.665 72.930 -86.480 ;
        RECT 73.505 -86.665 73.675 -86.650 ;
        RECT 66.100 -86.855 66.990 -86.685 ;
        RECT 72.760 -86.835 73.675 -86.665 ;
        RECT 66.100 -87.030 66.270 -86.855 ;
        RECT 65.155 -92.925 66.405 -92.350 ;
        RECT 66.810 -92.420 66.980 -86.855 ;
        RECT 72.760 -87.010 72.930 -86.835 ;
        RECT 66.730 -92.925 70.340 -92.895 ;
        RECT 65.155 -93.225 70.340 -92.925 ;
        RECT 71.885 -92.900 73.135 -92.350 ;
        RECT 73.505 -92.420 73.675 -86.835 ;
        RECT 78.875 -86.705 79.045 -86.520 ;
        RECT 79.620 -86.705 79.790 -86.650 ;
        RECT 78.875 -86.875 79.790 -86.705 ;
        RECT 78.875 -87.050 79.045 -86.875 ;
        RECT 77.980 -92.895 79.230 -92.350 ;
        RECT 79.620 -92.420 79.790 -86.875 ;
        RECT 85.300 -86.665 85.470 -86.480 ;
        RECT 86.025 -86.665 86.195 -86.650 ;
        RECT 85.300 -86.835 86.195 -86.665 ;
        RECT 85.300 -87.010 85.470 -86.835 ;
        RECT 73.425 -92.900 77.035 -92.895 ;
        RECT 71.885 -93.220 77.035 -92.900 ;
        RECT 65.155 -93.600 66.405 -93.225 ;
        RECT 71.885 -93.600 73.135 -93.220 ;
        RECT 73.425 -93.225 77.035 -93.220 ;
        RECT 77.980 -93.215 83.150 -92.895 ;
        RECT 77.980 -93.600 79.230 -93.215 ;
        RECT 79.540 -93.225 83.150 -93.215 ;
        RECT 84.350 -92.910 85.600 -92.180 ;
        RECT 86.025 -92.420 86.195 -86.835 ;
        RECT 85.945 -92.910 89.555 -92.895 ;
        RECT 84.350 -93.210 89.555 -92.910 ;
        RECT 84.350 -93.430 85.600 -93.210 ;
        RECT 85.945 -93.225 89.555 -93.210 ;
      LAYER met1 ;
        RECT 76.480 -59.200 77.120 -59.180 ;
        RECT 76.320 -60.100 77.280 -59.200 ;
        RECT 76.480 -60.120 77.120 -60.100 ;
        RECT 74.565 -72.280 75.205 -72.260 ;
        RECT 74.405 -73.180 75.365 -72.280 ;
        RECT 74.565 -73.200 75.205 -73.180 ;
        RECT 83.325 -73.320 83.975 -67.135 ;
        RECT 83.325 -73.970 93.975 -73.320 ;
        RECT 39.400 -78.405 40.040 -78.385 ;
        RECT 45.940 -78.405 46.580 -78.385 ;
        RECT 52.635 -78.405 53.275 -78.385 ;
        RECT 39.240 -79.305 40.200 -78.405 ;
        RECT 45.780 -79.305 46.740 -78.405 ;
        RECT 52.475 -79.305 53.435 -78.405 ;
        RECT 59.565 -78.480 60.205 -78.460 ;
        RECT 39.400 -79.325 40.040 -79.305 ;
        RECT 45.940 -79.325 46.580 -79.305 ;
        RECT 52.635 -79.325 53.275 -79.305 ;
        RECT 59.405 -79.380 60.365 -78.480 ;
        RECT 59.565 -79.400 60.205 -79.380 ;
        RECT 78.660 -80.550 79.300 -80.530 ;
        RECT 85.065 -80.550 85.705 -80.530 ;
        RECT 78.500 -81.450 79.460 -80.550 ;
        RECT 84.905 -81.450 85.865 -80.550 ;
        RECT 78.660 -81.470 79.300 -81.450 ;
        RECT 85.065 -81.470 85.705 -81.450 ;
        RECT 65.870 -81.740 66.510 -81.720 ;
        RECT 72.500 -81.740 73.140 -81.720 ;
        RECT 65.710 -82.640 66.670 -81.740 ;
        RECT 72.340 -82.640 73.300 -81.740 ;
        RECT 65.870 -82.660 66.510 -82.640 ;
        RECT 72.500 -82.660 73.140 -82.640 ;
        RECT 68.010 -83.240 68.650 -83.220 ;
        RECT 74.975 -83.240 75.615 -83.220 ;
        RECT 81.260 -83.240 81.900 -83.220 ;
        RECT 87.335 -83.240 87.975 -83.220 ;
        RECT 2.250 -84.090 2.890 -84.070 ;
        RECT 11.100 -84.090 11.740 -84.070 ;
        RECT 22.320 -84.090 22.960 -84.070 ;
        RECT 31.395 -84.090 32.035 -84.070 ;
        RECT 2.090 -84.990 3.050 -84.090 ;
        RECT 10.940 -84.990 11.900 -84.090 ;
        RECT 22.160 -84.990 23.120 -84.090 ;
        RECT 31.235 -84.990 32.195 -84.090 ;
        RECT 67.850 -84.140 68.810 -83.240 ;
        RECT 74.815 -84.140 75.775 -83.240 ;
        RECT 81.100 -84.140 82.060 -83.240 ;
        RECT 87.175 -84.140 88.135 -83.240 ;
        RECT 68.010 -84.160 68.650 -84.140 ;
        RECT 74.975 -84.160 75.615 -84.140 ;
        RECT 81.260 -84.160 81.900 -84.140 ;
        RECT 87.335 -84.160 87.975 -84.140 ;
        RECT 2.250 -85.010 2.890 -84.990 ;
        RECT 11.100 -85.010 11.740 -84.990 ;
        RECT 22.320 -85.010 22.960 -84.990 ;
        RECT 31.395 -85.010 32.035 -84.990 ;
        RECT 4.765 -85.845 5.405 -85.825 ;
        RECT 14.560 -85.845 15.200 -85.825 ;
        RECT 23.920 -85.845 24.560 -85.825 ;
        RECT 4.605 -86.745 5.565 -85.845 ;
        RECT 14.400 -86.745 15.360 -85.845 ;
        RECT 23.760 -86.745 24.720 -85.845 ;
        RECT 72.525 -86.295 73.165 -86.275 ;
        RECT 85.065 -86.295 85.705 -86.275 ;
        RECT 65.865 -86.315 66.505 -86.295 ;
        RECT 34.405 -86.450 35.045 -86.430 ;
        RECT 4.765 -86.765 5.405 -86.745 ;
        RECT 14.560 -86.765 15.200 -86.745 ;
        RECT 23.920 -86.765 24.560 -86.745 ;
        RECT 34.245 -87.350 35.205 -86.450 ;
        RECT 65.705 -87.215 66.665 -86.315 ;
        RECT 72.365 -87.195 73.325 -86.295 ;
        RECT 78.640 -86.335 79.280 -86.315 ;
        RECT 72.525 -87.215 73.165 -87.195 ;
        RECT 65.865 -87.235 66.505 -87.215 ;
        RECT 78.480 -87.235 79.440 -86.335 ;
        RECT 84.905 -87.195 85.865 -86.295 ;
        RECT 85.065 -87.215 85.705 -87.195 ;
        RECT 78.640 -87.255 79.280 -87.235 ;
        RECT 34.405 -87.370 35.045 -87.350 ;
        RECT 21.965 -93.665 22.605 -93.085 ;
        RECT 53.225 -93.150 53.865 -92.860 ;
        RECT 22.215 -94.145 22.355 -93.665 ;
        RECT 53.210 -94.145 53.910 -93.150 ;
        RECT 63.885 -94.145 64.585 -92.860 ;
        RECT 65.095 -93.630 66.465 -92.320 ;
        RECT 71.825 -93.630 73.195 -92.320 ;
        RECT 77.920 -93.630 79.290 -92.320 ;
        RECT 84.290 -93.460 85.660 -92.150 ;
        RECT 65.440 -94.145 66.140 -93.630 ;
        RECT 72.020 -94.145 72.720 -93.630 ;
        RECT 78.515 -94.145 79.215 -93.630 ;
        RECT 84.740 -94.145 85.440 -93.460 ;
        RECT 93.325 -94.145 93.975 -73.970 ;
        RECT 0.000 -100.255 99.790 -94.145 ;
      LAYER met2 ;
        RECT 76.320 -59.300 77.280 -59.200 ;
        RECT 73.425 -60.000 77.280 -59.300 ;
        RECT 73.425 -72.165 74.125 -60.000 ;
        RECT 76.320 -60.100 77.280 -60.000 ;
        RECT 73.425 -72.280 75.235 -72.165 ;
        RECT 73.425 -72.865 75.365 -72.280 ;
        RECT 74.405 -73.180 75.365 -72.865 ;
        RECT 74.535 -74.185 75.235 -73.180 ;
        RECT 65.825 -74.885 75.235 -74.185 ;
        RECT 39.240 -79.305 40.200 -78.405 ;
        RECT 45.780 -79.305 46.740 -78.405 ;
        RECT 52.475 -79.305 53.435 -78.405 ;
        RECT 39.260 -79.895 39.400 -79.305 ;
        RECT 45.825 -79.895 45.965 -79.305 ;
        RECT 52.545 -79.895 52.685 -79.305 ;
        RECT 59.405 -79.380 60.365 -78.480 ;
        RECT 59.435 -79.895 59.575 -79.380 ;
        RECT 39.260 -80.035 59.575 -79.895 ;
        RECT 2.090 -84.990 3.050 -84.090 ;
        RECT 10.940 -84.990 11.900 -84.090 ;
        RECT 22.160 -84.540 23.120 -84.090 ;
        RECT 21.975 -84.990 23.120 -84.540 ;
        RECT 31.235 -84.990 32.195 -84.090 ;
        RECT 2.280 -86.745 2.980 -84.990 ;
        RECT 10.955 -85.120 11.690 -84.990 ;
        RECT 4.605 -86.745 5.565 -85.845 ;
        RECT 10.955 -86.745 11.655 -85.120 ;
        RECT 14.400 -86.745 15.360 -85.845 ;
        RECT 21.975 -86.745 22.675 -84.990 ;
        RECT 23.760 -86.745 24.720 -85.845 ;
        RECT 31.405 -86.745 32.105 -84.990 ;
        RECT 34.245 -86.745 35.205 -86.450 ;
        RECT 2.280 -87.350 35.205 -86.745 ;
        RECT 2.280 -87.445 35.075 -87.350 ;
        RECT 21.975 -93.085 22.675 -87.445 ;
        RECT 21.965 -93.375 22.675 -93.085 ;
        RECT 21.965 -93.665 22.605 -93.375 ;
        RECT 53.195 -93.440 53.895 -80.035 ;
        RECT 65.825 -81.740 66.525 -74.885 ;
        RECT 78.500 -81.450 79.460 -80.550 ;
        RECT 84.905 -81.450 85.865 -80.550 ;
        RECT 65.710 -82.640 66.670 -81.740 ;
        RECT 72.340 -82.640 73.300 -81.740 ;
        RECT 65.840 -84.340 66.540 -82.640 ;
        RECT 67.850 -84.140 68.810 -83.240 ;
        RECT 68.180 -84.340 68.480 -84.140 ;
        RECT 72.670 -84.340 72.970 -82.640 ;
        RECT 74.815 -84.140 75.775 -83.240 ;
        RECT 75.145 -84.340 75.445 -84.140 ;
        RECT 79.190 -84.340 79.330 -81.450 ;
        RECT 81.100 -84.140 82.060 -83.240 ;
        RECT 85.300 -83.540 85.600 -81.450 ;
        RECT 87.175 -83.540 88.135 -83.240 ;
        RECT 85.300 -83.840 88.135 -83.540 ;
        RECT 81.430 -84.340 81.730 -84.140 ;
        RECT 85.300 -84.340 85.600 -83.840 ;
        RECT 87.175 -84.140 88.135 -83.840 ;
        RECT 65.840 -84.640 85.600 -84.340 ;
        RECT 65.840 -85.945 66.540 -84.640 ;
        RECT 65.840 -86.085 85.645 -85.945 ;
        RECT 65.840 -86.315 66.540 -86.085 ;
        RECT 72.695 -86.295 72.995 -86.085 ;
        RECT 65.705 -86.415 66.665 -86.315 ;
        RECT 63.965 -87.115 66.665 -86.415 ;
        RECT 63.965 -92.800 64.665 -87.115 ;
        RECT 65.705 -87.215 66.665 -87.115 ;
        RECT 72.365 -87.195 73.325 -86.295 ;
        RECT 79.015 -86.335 79.315 -86.085 ;
        RECT 85.505 -86.295 85.645 -86.085 ;
        RECT 78.480 -87.235 79.440 -86.335 ;
        RECT 84.905 -87.195 85.865 -86.295 ;
        RECT 63.915 -93.500 64.665 -92.800 ;
    END
  END Vss
  PIN Vout
    ANTENNADIFFAREA 17.639999 ;
    PORT
      LAYER li1 ;
        RECT 55.445 -18.230 55.615 -10.525 ;
        RECT 53.765 -18.300 55.615 -18.230 ;
        RECT 53.350 -18.400 55.615 -18.300 ;
        RECT 53.350 -19.300 54.350 -18.400 ;
        RECT 56.705 -19.180 56.875 -10.525 ;
        RECT 55.350 -19.350 56.875 -19.180 ;
        RECT 55.350 -20.360 55.520 -19.350 ;
        RECT 57.965 -20.155 58.135 -10.525 ;
        RECT 54.560 -20.530 55.520 -20.360 ;
        RECT 56.375 -20.325 58.135 -20.155 ;
        RECT 53.350 -21.395 54.350 -21.300 ;
        RECT 54.560 -21.395 54.730 -20.530 ;
        RECT 56.375 -21.380 56.545 -20.325 ;
        RECT 59.225 -21.250 59.395 -10.525 ;
        RECT 53.350 -21.565 54.730 -21.395 ;
        RECT 55.755 -21.550 56.545 -21.380 ;
        RECT 57.780 -21.420 59.395 -21.250 ;
        RECT 53.350 -22.300 54.350 -21.565 ;
        RECT 55.755 -22.410 55.925 -21.550 ;
        RECT 55.230 -22.580 55.925 -22.410 ;
        RECT 55.230 -23.550 55.400 -22.580 ;
        RECT 54.760 -24.550 55.760 -23.550 ;
        RECT 56.435 -24.045 57.435 -23.885 ;
        RECT 57.780 -24.045 57.950 -21.420 ;
        RECT 60.485 -23.885 60.655 -10.525 ;
        RECT 61.745 -17.150 61.915 -10.525 ;
        RECT 61.735 -17.315 61.915 -17.150 ;
        RECT 61.735 -21.370 61.905 -17.315 ;
        RECT 63.005 -20.235 63.175 -10.525 ;
        RECT 64.265 -19.160 64.435 -10.525 ;
        RECT 65.525 -17.940 65.695 -10.525 ;
        RECT 65.525 -18.070 67.430 -17.940 ;
        RECT 65.525 -18.110 67.860 -18.070 ;
        RECT 66.860 -19.070 67.860 -18.110 ;
        RECT 64.265 -19.330 65.700 -19.160 ;
        RECT 65.530 -19.955 65.700 -19.330 ;
        RECT 65.530 -20.125 66.575 -19.955 ;
        RECT 63.005 -20.405 64.510 -20.235 ;
        RECT 64.340 -21.015 64.510 -20.405 ;
        RECT 66.405 -20.790 66.575 -20.125 ;
        RECT 66.405 -20.800 67.485 -20.790 ;
        RECT 66.405 -20.960 67.900 -20.800 ;
        RECT 64.340 -21.185 65.510 -21.015 ;
        RECT 61.735 -21.540 63.215 -21.370 ;
        RECT 63.045 -22.165 63.215 -21.540 ;
        RECT 65.340 -22.005 65.510 -21.185 ;
        RECT 66.900 -21.800 67.900 -20.960 ;
        RECT 63.045 -22.335 63.470 -22.165 ;
        RECT 65.340 -22.175 66.065 -22.005 ;
        RECT 56.435 -24.215 57.950 -24.045 ;
        RECT 56.435 -24.885 57.435 -24.215 ;
        RECT 60.055 -24.885 61.055 -23.885 ;
        RECT 63.300 -24.300 63.470 -22.335 ;
        RECT 65.895 -23.210 66.065 -22.175 ;
        RECT 63.805 -24.300 64.805 -23.885 ;
        RECT 65.410 -24.210 66.410 -23.210 ;
        RECT 63.300 -24.470 64.805 -24.300 ;
        RECT 63.805 -24.885 64.805 -24.470 ;
        RECT 88.155 -42.270 88.825 -42.100 ;
      LAYER met1 ;
        RECT 53.350 -19.300 54.350 -18.300 ;
        RECT 66.860 -19.070 67.860 -18.070 ;
        RECT 53.350 -22.300 54.350 -21.300 ;
        RECT 66.900 -21.800 67.900 -20.800 ;
        RECT 54.760 -24.550 55.760 -23.550 ;
        RECT 56.435 -24.885 57.435 -23.885 ;
        RECT 60.055 -24.885 61.055 -23.885 ;
        RECT 63.805 -24.885 64.805 -23.885 ;
        RECT 65.410 -24.210 66.410 -23.210 ;
        RECT 91.780 -33.675 92.780 -32.675 ;
        RECT 91.955 -41.090 92.605 -33.675 ;
        RECT 94.540 -41.090 99.780 -32.620 ;
        RECT 88.165 -41.740 99.780 -41.090 ;
        RECT 88.165 -42.300 88.815 -41.740 ;
        RECT 94.540 -42.620 99.780 -41.740 ;
      LAYER met2 ;
        RECT 53.265 -19.365 54.435 -18.235 ;
        RECT 66.775 -19.135 67.945 -18.005 ;
        RECT 53.265 -22.365 54.435 -21.235 ;
        RECT 66.815 -21.865 67.985 -20.735 ;
        RECT 54.675 -24.615 55.845 -23.485 ;
        RECT 56.350 -24.950 57.520 -23.820 ;
        RECT 59.970 -24.950 61.140 -23.820 ;
        RECT 63.720 -24.950 64.890 -23.820 ;
        RECT 65.325 -24.275 66.495 -23.145 ;
        RECT 91.695 -33.740 92.865 -32.610 ;
      LAYER met3 ;
        RECT 66.775 -18.235 67.945 -18.005 ;
        RECT 53.265 -18.450 54.435 -18.235 ;
        RECT 51.480 -19.150 54.435 -18.450 ;
        RECT 66.775 -18.935 70.235 -18.235 ;
        RECT 66.775 -19.135 67.945 -18.935 ;
        RECT 51.480 -21.050 52.180 -19.150 ;
        RECT 53.265 -19.365 54.435 -19.150 ;
        RECT 51.450 -21.430 52.180 -21.050 ;
        RECT 66.815 -20.950 67.985 -20.735 ;
        RECT 69.535 -20.950 70.235 -18.935 ;
        RECT 53.265 -21.430 54.435 -21.235 ;
        RECT 51.450 -22.130 54.435 -21.430 ;
        RECT 66.815 -21.650 70.235 -20.950 ;
        RECT 66.815 -21.865 67.985 -21.650 ;
        RECT 51.450 -25.020 52.150 -22.130 ;
        RECT 53.265 -22.365 54.435 -22.130 ;
        RECT 54.675 -24.615 55.845 -23.485 ;
        RECT 54.895 -25.020 55.595 -24.615 ;
        RECT 56.350 -24.950 57.520 -23.820 ;
        RECT 59.970 -24.950 61.140 -23.820 ;
        RECT 63.720 -24.595 64.890 -23.820 ;
        RECT 65.325 -24.275 66.495 -23.145 ;
        RECT 65.560 -24.595 66.260 -24.275 ;
        RECT 68.645 -24.595 68.945 -24.455 ;
        RECT 63.720 -24.655 68.945 -24.595 ;
        RECT 69.535 -24.655 70.235 -21.650 ;
        RECT 63.720 -24.950 70.235 -24.655 ;
        RECT 51.450 -25.720 55.595 -25.020 ;
        RECT 54.895 -26.215 55.595 -25.720 ;
        RECT 56.785 -26.215 57.085 -24.950 ;
        RECT 60.405 -26.150 60.705 -24.950 ;
        RECT 63.955 -24.955 70.235 -24.950 ;
        RECT 63.955 -25.295 68.945 -24.955 ;
        RECT 59.825 -26.155 60.705 -26.150 ;
        RECT 65.560 -26.155 66.260 -25.295 ;
        RECT 59.825 -26.215 66.260 -26.155 ;
        RECT 54.895 -26.855 66.260 -26.215 ;
        RECT 54.895 -26.915 60.525 -26.855 ;
        RECT 69.535 -32.930 70.235 -24.955 ;
        RECT 91.695 -32.930 92.865 -32.610 ;
        RECT 69.535 -33.630 92.865 -32.930 ;
        RECT 91.695 -33.740 92.865 -33.630 ;
    END
  END Vout
  PIN Vinp
    ANTENNAGATEAREA 4.410000 ;
    PORT
      LAYER li1 ;
        RECT 76.510 -50.240 77.180 -49.630 ;
      LAYER met1 ;
        RECT 94.710 -49.595 99.785 -49.585 ;
        RECT 76.450 -50.295 99.785 -49.595 ;
        RECT 94.710 -59.585 99.785 -50.295 ;
    END
  END Vinp
  PIN Vinn
    ANTENNAGATEAREA 4.410000 ;
    PORT
      LAYER li1 ;
        RECT 76.630 -64.290 77.300 -63.680 ;
      LAYER met1 ;
        RECT 94.525 -63.550 99.805 -63.525 ;
        RECT 76.700 -63.690 99.805 -63.550 ;
        RECT 76.640 -64.250 99.805 -63.690 ;
        RECT 76.640 -64.280 77.290 -64.250 ;
        RECT 94.525 -73.525 99.805 -64.250 ;
    END
  END Vinn
  OBS
      LAYER li1 ;
        RECT 6.470 -7.055 8.350 -6.885 ;
        RECT 8.890 -7.055 10.770 -6.885 ;
        RECT 15.545 -14.025 15.715 -13.845 ;
        RECT 16.620 -14.025 16.790 -9.735 ;
        RECT 15.545 -14.195 16.790 -14.025 ;
        RECT 15.545 -14.375 15.715 -14.195 ;
        RECT 16.620 -14.485 16.790 -14.195 ;
        RECT 17.250 -14.370 17.420 -9.735 ;
        RECT 17.250 -14.485 17.430 -14.370 ;
        RECT 14.935 -15.170 15.935 -15.065 ;
        RECT 17.260 -15.170 17.430 -14.485 ;
        RECT 14.935 -15.340 17.430 -15.170 ;
        RECT 14.935 -16.065 15.935 -15.340 ;
        RECT 17.880 -15.690 18.050 -9.735 ;
        RECT 18.510 -14.800 18.680 -9.735 ;
        RECT 19.140 -14.785 19.310 -9.735 ;
        RECT 16.820 -15.775 18.050 -15.690 ;
        RECT 16.795 -15.860 18.050 -15.775 ;
        RECT 18.295 -14.970 18.680 -14.800 ;
        RECT 18.940 -14.955 19.310 -14.785 ;
        RECT 16.795 -15.935 16.990 -15.860 ;
        RECT 16.795 -16.305 16.965 -15.935 ;
        RECT 18.295 -16.130 18.465 -14.970 ;
        RECT 18.940 -15.260 19.110 -14.955 ;
        RECT 17.635 -16.300 18.465 -16.130 ;
        RECT 18.700 -15.430 19.110 -15.260 ;
        RECT 19.770 -15.365 19.940 -9.735 ;
        RECT 17.635 -16.970 17.805 -16.300 ;
        RECT 18.700 -16.740 18.870 -15.430 ;
        RECT 16.660 -17.395 17.805 -16.970 ;
        RECT 18.465 -16.910 18.870 -16.740 ;
        RECT 19.330 -15.535 19.940 -15.365 ;
        RECT 18.465 -17.355 18.635 -16.910 ;
        RECT 16.660 -17.970 17.660 -17.395 ;
        RECT 19.330 -18.000 19.500 -15.535 ;
        RECT 20.400 -15.725 20.570 -9.735 ;
        RECT 14.745 -18.565 15.275 -18.035 ;
        RECT 18.225 -18.170 19.500 -18.000 ;
        RECT 19.810 -15.895 20.570 -15.725 ;
        RECT 18.225 -19.000 19.225 -18.170 ;
        RECT 19.810 -18.940 19.980 -15.895 ;
        RECT 21.030 -16.450 21.200 -9.735 ;
        RECT 20.335 -16.620 21.200 -16.450 ;
        RECT 20.335 -18.145 20.505 -16.620 ;
        RECT 20.335 -18.315 21.225 -18.145 ;
        RECT 19.810 -19.110 20.215 -18.940 ;
        RECT 20.045 -19.470 20.215 -19.110 ;
        RECT 19.730 -20.530 20.730 -20.350 ;
        RECT 21.055 -20.530 21.225 -18.315 ;
        RECT 21.660 -18.785 21.830 -9.735 ;
        RECT 19.730 -20.700 21.225 -20.530 ;
        RECT 21.490 -18.955 21.830 -18.785 ;
        RECT 19.730 -21.350 20.730 -20.700 ;
        RECT 21.490 -20.890 21.660 -18.955 ;
        RECT 21.490 -21.060 21.685 -20.890 ;
        RECT 21.515 -21.880 21.685 -21.060 ;
        RECT 20.945 -22.050 21.685 -21.880 ;
        RECT 20.945 -22.140 21.115 -22.050 ;
        RECT 20.860 -22.670 21.115 -22.140 ;
        RECT 22.290 -23.565 22.460 -9.735 ;
        RECT 22.920 -14.285 23.090 -9.735 ;
        RECT 22.920 -14.485 23.120 -14.285 ;
        RECT 23.550 -14.335 23.720 -9.735 ;
        RECT 22.950 -15.870 23.120 -14.485 ;
        RECT 23.535 -14.485 23.720 -14.335 ;
        RECT 24.180 -14.345 24.350 -9.735 ;
        RECT 24.180 -14.485 24.370 -14.345 ;
        RECT 23.535 -15.305 23.705 -14.485 ;
        RECT 24.200 -14.845 24.370 -14.485 ;
        RECT 24.200 -15.015 24.410 -14.845 ;
        RECT 23.535 -15.475 23.925 -15.305 ;
        RECT 22.950 -16.040 23.390 -15.870 ;
        RECT 23.220 -22.670 23.390 -16.040 ;
        RECT 23.755 -21.445 23.925 -15.475 ;
        RECT 24.240 -19.720 24.410 -15.015 ;
        RECT 24.810 -19.065 24.980 -9.735 ;
        RECT 25.440 -17.600 25.610 -9.735 ;
        RECT 26.070 -16.890 26.240 -9.735 ;
        RECT 26.700 -16.280 26.870 -9.735 ;
        RECT 27.330 -15.660 27.500 -9.735 ;
        RECT 27.960 -15.170 28.130 -9.735 ;
        RECT 28.590 -13.945 28.760 -9.735 ;
        RECT 29.180 -13.945 30.180 -13.530 ;
        RECT 28.590 -14.115 30.180 -13.945 ;
        RECT 28.590 -14.485 28.760 -14.115 ;
        RECT 29.180 -14.530 30.180 -14.115 ;
        RECT 34.080 -13.995 34.250 -13.815 ;
        RECT 35.155 -13.995 35.325 -9.730 ;
        RECT 34.080 -14.165 35.325 -13.995 ;
        RECT 34.080 -14.345 34.250 -14.165 ;
        RECT 35.155 -14.480 35.325 -14.165 ;
        RECT 35.785 -14.340 35.955 -9.730 ;
        RECT 35.785 -14.480 35.965 -14.340 ;
        RECT 33.470 -15.140 34.470 -15.035 ;
        RECT 35.795 -15.140 35.965 -14.480 ;
        RECT 27.960 -15.340 29.625 -15.170 ;
        RECT 29.455 -15.415 29.625 -15.340 ;
        RECT 33.470 -15.310 35.965 -15.140 ;
        RECT 27.330 -15.830 28.685 -15.660 ;
        RECT 29.455 -15.765 29.660 -15.415 ;
        RECT 26.700 -16.450 28.130 -16.280 ;
        RECT 26.070 -17.060 27.280 -16.890 ;
        RECT 25.440 -17.770 26.415 -17.600 ;
        RECT 26.205 -18.050 26.415 -17.770 ;
        RECT 26.205 -18.230 26.375 -18.050 ;
        RECT 27.110 -18.910 27.280 -17.060 ;
        RECT 27.960 -17.495 28.130 -16.450 ;
        RECT 28.515 -16.720 28.685 -15.830 ;
        RECT 29.490 -15.945 29.660 -15.765 ;
        RECT 33.470 -16.035 34.470 -15.310 ;
        RECT 36.415 -15.660 36.585 -9.730 ;
        RECT 37.045 -14.770 37.215 -9.730 ;
        RECT 37.675 -14.755 37.845 -9.730 ;
        RECT 35.355 -15.745 36.585 -15.660 ;
        RECT 35.330 -15.830 36.585 -15.745 ;
        RECT 36.830 -14.940 37.215 -14.770 ;
        RECT 37.475 -14.925 37.845 -14.755 ;
        RECT 35.330 -15.905 35.525 -15.830 ;
        RECT 35.330 -16.275 35.500 -15.905 ;
        RECT 36.830 -16.100 37.000 -14.940 ;
        RECT 37.475 -15.230 37.645 -14.925 ;
        RECT 36.170 -16.270 37.000 -16.100 ;
        RECT 37.235 -15.400 37.645 -15.230 ;
        RECT 38.305 -15.335 38.475 -9.730 ;
        RECT 29.180 -16.720 30.180 -16.685 ;
        RECT 28.515 -16.890 30.180 -16.720 ;
        RECT 27.960 -17.845 28.200 -17.495 ;
        RECT 29.180 -17.685 30.180 -16.890 ;
        RECT 36.170 -16.940 36.340 -16.270 ;
        RECT 37.235 -16.710 37.405 -15.400 ;
        RECT 35.195 -17.365 36.340 -16.940 ;
        RECT 37.000 -16.880 37.405 -16.710 ;
        RECT 37.865 -15.505 38.475 -15.335 ;
        RECT 37.000 -17.325 37.170 -16.880 ;
        RECT 28.030 -18.025 28.200 -17.845 ;
        RECT 35.195 -17.940 36.195 -17.365 ;
        RECT 37.865 -17.970 38.035 -15.505 ;
        RECT 38.935 -15.695 39.105 -9.730 ;
        RECT 36.760 -18.140 38.035 -17.970 ;
        RECT 38.345 -15.865 39.105 -15.695 ;
        RECT 27.110 -18.955 28.225 -18.910 ;
        RECT 25.695 -19.065 26.695 -18.955 ;
        RECT 24.810 -19.235 26.695 -19.065 ;
        RECT 27.110 -19.080 28.640 -18.955 ;
        RECT 24.240 -19.890 24.855 -19.720 ;
        RECT 24.685 -20.335 24.855 -19.890 ;
        RECT 25.695 -19.955 26.695 -19.235 ;
        RECT 27.640 -19.955 28.640 -19.080 ;
        RECT 34.100 -19.260 34.630 -18.730 ;
        RECT 36.760 -18.970 37.760 -18.140 ;
        RECT 38.345 -18.910 38.515 -15.865 ;
        RECT 39.565 -16.420 39.735 -9.730 ;
        RECT 38.870 -16.590 39.735 -16.420 ;
        RECT 38.870 -18.115 39.040 -16.590 ;
        RECT 38.870 -18.285 39.760 -18.115 ;
        RECT 38.345 -19.080 38.750 -18.910 ;
        RECT 38.580 -19.440 38.750 -19.080 ;
        RECT 38.265 -20.500 39.265 -20.320 ;
        RECT 39.590 -20.500 39.760 -18.285 ;
        RECT 40.195 -18.755 40.365 -9.730 ;
        RECT 38.265 -20.670 39.760 -20.500 ;
        RECT 40.025 -18.925 40.365 -18.755 ;
        RECT 24.270 -21.445 25.270 -21.030 ;
        RECT 38.265 -21.320 39.265 -20.670 ;
        RECT 40.025 -20.860 40.195 -18.925 ;
        RECT 40.025 -21.030 40.220 -20.860 ;
        RECT 23.755 -21.615 25.270 -21.445 ;
        RECT 24.270 -22.030 25.270 -21.615 ;
        RECT 40.050 -21.850 40.220 -21.030 ;
        RECT 39.480 -22.020 40.220 -21.850 ;
        RECT 39.480 -22.110 39.650 -22.020 ;
        RECT 39.395 -22.640 39.650 -22.110 ;
        RECT 40.825 -23.535 40.995 -9.730 ;
        RECT 41.455 -14.255 41.625 -9.730 ;
        RECT 41.455 -14.480 41.655 -14.255 ;
        RECT 42.085 -14.305 42.255 -9.730 ;
        RECT 41.485 -15.840 41.655 -14.480 ;
        RECT 42.070 -14.480 42.255 -14.305 ;
        RECT 42.715 -14.315 42.885 -9.730 ;
        RECT 42.715 -14.480 42.905 -14.315 ;
        RECT 42.070 -15.275 42.240 -14.480 ;
        RECT 42.735 -14.815 42.905 -14.480 ;
        RECT 42.735 -14.985 42.945 -14.815 ;
        RECT 42.070 -15.445 42.460 -15.275 ;
        RECT 41.485 -16.010 41.925 -15.840 ;
        RECT 41.755 -22.640 41.925 -16.010 ;
        RECT 42.290 -21.415 42.460 -15.445 ;
        RECT 42.775 -19.690 42.945 -14.985 ;
        RECT 43.345 -19.035 43.515 -9.730 ;
        RECT 43.975 -17.570 44.145 -9.730 ;
        RECT 44.605 -16.860 44.775 -9.730 ;
        RECT 45.235 -16.250 45.405 -9.730 ;
        RECT 45.865 -15.630 46.035 -9.730 ;
        RECT 46.495 -15.140 46.665 -9.730 ;
        RECT 47.125 -13.915 47.295 -9.730 ;
        RECT 47.715 -13.915 48.715 -13.500 ;
        RECT 47.125 -14.085 48.715 -13.915 ;
        RECT 47.125 -14.480 47.295 -14.085 ;
        RECT 47.715 -14.500 48.715 -14.085 ;
        RECT 46.495 -15.310 48.160 -15.140 ;
        RECT 47.990 -15.385 48.160 -15.310 ;
        RECT 45.865 -15.800 47.220 -15.630 ;
        RECT 47.990 -15.735 48.195 -15.385 ;
        RECT 45.235 -16.420 46.665 -16.250 ;
        RECT 44.605 -17.030 45.815 -16.860 ;
        RECT 43.975 -17.740 44.950 -17.570 ;
        RECT 44.740 -18.020 44.950 -17.740 ;
        RECT 44.740 -18.200 44.910 -18.020 ;
        RECT 45.645 -18.880 45.815 -17.030 ;
        RECT 46.495 -17.465 46.665 -16.420 ;
        RECT 47.050 -16.690 47.220 -15.800 ;
        RECT 48.025 -15.915 48.195 -15.735 ;
        RECT 47.715 -16.690 48.715 -16.655 ;
        RECT 47.050 -16.860 48.715 -16.690 ;
        RECT 46.495 -17.815 46.735 -17.465 ;
        RECT 47.715 -17.655 48.715 -16.860 ;
        RECT 46.565 -17.995 46.735 -17.815 ;
        RECT 69.360 -18.085 69.890 -17.555 ;
        RECT 45.645 -18.925 46.760 -18.880 ;
        RECT 44.230 -19.035 45.230 -18.925 ;
        RECT 43.345 -19.205 45.230 -19.035 ;
        RECT 45.645 -19.050 47.175 -18.925 ;
        RECT 42.775 -19.860 43.390 -19.690 ;
        RECT 43.220 -20.305 43.390 -19.860 ;
        RECT 44.230 -19.925 45.230 -19.205 ;
        RECT 46.175 -19.925 47.175 -19.050 ;
        RECT 42.805 -21.415 43.805 -21.000 ;
        RECT 42.290 -21.585 43.805 -21.415 ;
        RECT 42.805 -22.000 43.805 -21.585 ;
        RECT 21.870 -24.565 22.870 -23.565 ;
        RECT 40.390 -24.535 41.390 -23.535 ;
        RECT 15.545 -32.355 15.715 -32.175 ;
        RECT 16.620 -32.355 16.790 -28.080 ;
        RECT 15.545 -32.525 16.790 -32.355 ;
        RECT 15.545 -32.705 15.715 -32.525 ;
        RECT 16.620 -32.830 16.790 -32.525 ;
        RECT 17.250 -32.700 17.420 -28.080 ;
        RECT 17.250 -32.830 17.430 -32.700 ;
        RECT 14.935 -33.500 15.935 -33.395 ;
        RECT 17.260 -33.500 17.430 -32.830 ;
        RECT 14.935 -33.670 17.430 -33.500 ;
        RECT 14.935 -34.395 15.935 -33.670 ;
        RECT 17.880 -34.020 18.050 -28.080 ;
        RECT 18.510 -33.130 18.680 -28.080 ;
        RECT 19.140 -33.115 19.310 -28.080 ;
        RECT 16.820 -34.105 18.050 -34.020 ;
        RECT 16.795 -34.190 18.050 -34.105 ;
        RECT 18.295 -33.300 18.680 -33.130 ;
        RECT 18.940 -33.285 19.310 -33.115 ;
        RECT 16.795 -34.265 16.990 -34.190 ;
        RECT 16.795 -34.635 16.965 -34.265 ;
        RECT 18.295 -34.460 18.465 -33.300 ;
        RECT 18.940 -33.590 19.110 -33.285 ;
        RECT 17.635 -34.630 18.465 -34.460 ;
        RECT 18.700 -33.760 19.110 -33.590 ;
        RECT 19.770 -33.695 19.940 -28.080 ;
        RECT 17.635 -35.300 17.805 -34.630 ;
        RECT 18.700 -35.070 18.870 -33.760 ;
        RECT 16.660 -35.725 17.805 -35.300 ;
        RECT 18.465 -35.240 18.870 -35.070 ;
        RECT 19.330 -33.865 19.940 -33.695 ;
        RECT 18.465 -35.685 18.635 -35.240 ;
        RECT 16.660 -36.300 17.660 -35.725 ;
        RECT 19.330 -36.330 19.500 -33.865 ;
        RECT 20.400 -34.055 20.570 -28.080 ;
        RECT 18.225 -36.500 19.500 -36.330 ;
        RECT 19.810 -34.225 20.570 -34.055 ;
        RECT 15.340 -37.600 15.870 -37.070 ;
        RECT 18.225 -37.330 19.225 -36.500 ;
        RECT 19.810 -37.270 19.980 -34.225 ;
        RECT 21.030 -34.780 21.200 -28.080 ;
        RECT 20.335 -34.950 21.200 -34.780 ;
        RECT 20.335 -36.475 20.505 -34.950 ;
        RECT 20.335 -36.645 21.225 -36.475 ;
        RECT 19.810 -37.440 20.215 -37.270 ;
        RECT 20.045 -37.800 20.215 -37.440 ;
        RECT 19.730 -38.860 20.730 -38.680 ;
        RECT 21.055 -38.860 21.225 -36.645 ;
        RECT 21.660 -37.115 21.830 -28.080 ;
        RECT 19.730 -39.030 21.225 -38.860 ;
        RECT 21.490 -37.285 21.830 -37.115 ;
        RECT 19.730 -39.680 20.730 -39.030 ;
        RECT 21.490 -39.220 21.660 -37.285 ;
        RECT 21.490 -39.390 21.685 -39.220 ;
        RECT 21.515 -40.210 21.685 -39.390 ;
        RECT 20.945 -40.380 21.685 -40.210 ;
        RECT 20.945 -40.470 21.115 -40.380 ;
        RECT 20.860 -41.000 21.115 -40.470 ;
        RECT 22.290 -41.895 22.460 -28.080 ;
        RECT 22.920 -32.615 23.090 -28.080 ;
        RECT 22.920 -32.830 23.120 -32.615 ;
        RECT 23.550 -32.665 23.720 -28.080 ;
        RECT 22.950 -34.200 23.120 -32.830 ;
        RECT 23.535 -32.830 23.720 -32.665 ;
        RECT 24.180 -32.675 24.350 -28.080 ;
        RECT 24.180 -32.830 24.370 -32.675 ;
        RECT 23.535 -33.635 23.705 -32.830 ;
        RECT 24.200 -33.175 24.370 -32.830 ;
        RECT 24.200 -33.345 24.410 -33.175 ;
        RECT 23.535 -33.805 23.925 -33.635 ;
        RECT 22.950 -34.370 23.390 -34.200 ;
        RECT 23.220 -41.000 23.390 -34.370 ;
        RECT 23.755 -39.775 23.925 -33.805 ;
        RECT 24.240 -38.050 24.410 -33.345 ;
        RECT 24.810 -37.395 24.980 -28.080 ;
        RECT 25.440 -35.930 25.610 -28.080 ;
        RECT 26.070 -35.220 26.240 -28.080 ;
        RECT 26.700 -34.610 26.870 -28.080 ;
        RECT 27.330 -33.990 27.500 -28.080 ;
        RECT 27.960 -33.500 28.130 -28.080 ;
        RECT 28.590 -32.275 28.760 -28.080 ;
        RECT 29.180 -32.275 30.180 -31.860 ;
        RECT 28.590 -32.445 30.180 -32.275 ;
        RECT 28.590 -32.830 28.760 -32.445 ;
        RECT 29.180 -32.860 30.180 -32.445 ;
        RECT 33.835 -32.645 34.005 -32.465 ;
        RECT 34.910 -32.645 35.080 -28.385 ;
        RECT 33.835 -32.815 35.080 -32.645 ;
        RECT 33.835 -32.995 34.005 -32.815 ;
        RECT 34.910 -33.135 35.080 -32.815 ;
        RECT 35.540 -32.990 35.710 -28.385 ;
        RECT 35.540 -33.135 35.720 -32.990 ;
        RECT 27.960 -33.670 29.625 -33.500 ;
        RECT 29.455 -33.745 29.625 -33.670 ;
        RECT 27.330 -34.160 28.685 -33.990 ;
        RECT 29.455 -34.095 29.660 -33.745 ;
        RECT 26.700 -34.780 28.130 -34.610 ;
        RECT 26.070 -35.390 27.280 -35.220 ;
        RECT 25.440 -36.100 26.415 -35.930 ;
        RECT 26.205 -36.380 26.415 -36.100 ;
        RECT 26.205 -36.560 26.375 -36.380 ;
        RECT 27.110 -37.240 27.280 -35.390 ;
        RECT 27.960 -35.825 28.130 -34.780 ;
        RECT 28.515 -35.050 28.685 -34.160 ;
        RECT 29.490 -34.275 29.660 -34.095 ;
        RECT 33.225 -33.790 34.225 -33.635 ;
        RECT 35.550 -33.790 35.720 -33.135 ;
        RECT 33.225 -33.960 35.720 -33.790 ;
        RECT 33.225 -34.635 34.225 -33.960 ;
        RECT 36.170 -34.310 36.340 -28.385 ;
        RECT 36.800 -33.420 36.970 -28.385 ;
        RECT 37.430 -33.405 37.600 -28.385 ;
        RECT 35.110 -34.395 36.340 -34.310 ;
        RECT 35.085 -34.480 36.340 -34.395 ;
        RECT 36.585 -33.590 36.970 -33.420 ;
        RECT 37.230 -33.575 37.600 -33.405 ;
        RECT 35.085 -34.555 35.280 -34.480 ;
        RECT 35.085 -34.925 35.255 -34.555 ;
        RECT 36.585 -34.750 36.755 -33.590 ;
        RECT 37.230 -33.880 37.400 -33.575 ;
        RECT 35.925 -34.920 36.755 -34.750 ;
        RECT 36.990 -34.050 37.400 -33.880 ;
        RECT 38.060 -33.985 38.230 -28.385 ;
        RECT 29.180 -35.050 30.180 -35.015 ;
        RECT 28.515 -35.220 30.180 -35.050 ;
        RECT 27.960 -36.175 28.200 -35.825 ;
        RECT 29.180 -36.015 30.180 -35.220 ;
        RECT 35.925 -35.590 36.095 -34.920 ;
        RECT 36.990 -35.360 37.160 -34.050 ;
        RECT 34.950 -36.015 36.095 -35.590 ;
        RECT 36.755 -35.530 37.160 -35.360 ;
        RECT 37.620 -34.155 38.230 -33.985 ;
        RECT 36.755 -35.975 36.925 -35.530 ;
        RECT 28.030 -36.355 28.200 -36.175 ;
        RECT 34.950 -36.590 35.950 -36.015 ;
        RECT 37.620 -36.620 37.790 -34.155 ;
        RECT 38.690 -34.345 38.860 -28.385 ;
        RECT 36.515 -36.790 37.790 -36.620 ;
        RECT 38.100 -34.515 38.860 -34.345 ;
        RECT 27.110 -37.285 28.225 -37.240 ;
        RECT 25.695 -37.395 26.695 -37.285 ;
        RECT 24.810 -37.565 26.695 -37.395 ;
        RECT 27.110 -37.410 28.640 -37.285 ;
        RECT 24.240 -38.220 24.855 -38.050 ;
        RECT 24.685 -38.665 24.855 -38.220 ;
        RECT 25.695 -38.285 26.695 -37.565 ;
        RECT 27.640 -38.285 28.640 -37.410 ;
        RECT 33.725 -37.910 34.255 -37.380 ;
        RECT 36.515 -37.620 37.515 -36.790 ;
        RECT 38.100 -37.560 38.270 -34.515 ;
        RECT 39.320 -35.070 39.490 -28.385 ;
        RECT 38.625 -35.240 39.490 -35.070 ;
        RECT 38.625 -36.765 38.795 -35.240 ;
        RECT 38.625 -36.935 39.515 -36.765 ;
        RECT 38.100 -37.730 38.505 -37.560 ;
        RECT 38.335 -38.090 38.505 -37.730 ;
        RECT 38.020 -39.150 39.020 -38.970 ;
        RECT 39.345 -39.150 39.515 -36.935 ;
        RECT 39.950 -37.405 40.120 -28.385 ;
        RECT 38.020 -39.320 39.515 -39.150 ;
        RECT 39.780 -37.575 40.120 -37.405 ;
        RECT 24.270 -39.775 25.270 -39.360 ;
        RECT 23.755 -39.945 25.270 -39.775 ;
        RECT 24.270 -40.360 25.270 -39.945 ;
        RECT 38.020 -39.970 39.020 -39.320 ;
        RECT 39.780 -39.510 39.950 -37.575 ;
        RECT 39.780 -39.680 39.975 -39.510 ;
        RECT 39.805 -40.500 39.975 -39.680 ;
        RECT 39.235 -40.670 39.975 -40.500 ;
        RECT 39.235 -40.760 39.405 -40.670 ;
        RECT 39.150 -41.290 39.405 -40.760 ;
        RECT 21.890 -42.895 22.890 -41.895 ;
        RECT 40.580 -42.185 40.750 -28.385 ;
        RECT 41.210 -32.905 41.380 -28.385 ;
        RECT 41.210 -33.135 41.410 -32.905 ;
        RECT 41.840 -32.955 42.010 -28.385 ;
        RECT 41.240 -34.490 41.410 -33.135 ;
        RECT 41.825 -33.135 42.010 -32.955 ;
        RECT 42.470 -32.965 42.640 -28.385 ;
        RECT 42.470 -33.135 42.660 -32.965 ;
        RECT 41.825 -33.925 41.995 -33.135 ;
        RECT 42.490 -33.465 42.660 -33.135 ;
        RECT 42.490 -33.635 42.700 -33.465 ;
        RECT 41.825 -34.095 42.215 -33.925 ;
        RECT 41.240 -34.660 41.680 -34.490 ;
        RECT 41.510 -41.290 41.680 -34.660 ;
        RECT 42.045 -40.065 42.215 -34.095 ;
        RECT 42.530 -38.340 42.700 -33.635 ;
        RECT 43.100 -37.685 43.270 -28.385 ;
        RECT 43.730 -36.220 43.900 -28.385 ;
        RECT 44.360 -35.510 44.530 -28.385 ;
        RECT 44.990 -34.900 45.160 -28.385 ;
        RECT 45.620 -34.280 45.790 -28.385 ;
        RECT 46.250 -33.790 46.420 -28.385 ;
        RECT 46.880 -32.565 47.050 -28.385 ;
        RECT 47.470 -32.565 48.470 -32.150 ;
        RECT 46.880 -32.735 48.470 -32.565 ;
        RECT 46.880 -33.135 47.050 -32.735 ;
        RECT 47.470 -33.150 48.470 -32.735 ;
        RECT 46.250 -33.960 47.915 -33.790 ;
        RECT 47.745 -34.035 47.915 -33.960 ;
        RECT 45.620 -34.450 46.975 -34.280 ;
        RECT 47.745 -34.385 47.950 -34.035 ;
        RECT 44.990 -35.070 46.420 -34.900 ;
        RECT 44.360 -35.680 45.570 -35.510 ;
        RECT 43.730 -36.390 44.705 -36.220 ;
        RECT 44.495 -36.670 44.705 -36.390 ;
        RECT 44.495 -36.850 44.665 -36.670 ;
        RECT 45.400 -37.530 45.570 -35.680 ;
        RECT 46.250 -36.115 46.420 -35.070 ;
        RECT 46.805 -35.340 46.975 -34.450 ;
        RECT 47.780 -34.565 47.950 -34.385 ;
        RECT 47.470 -35.340 48.470 -35.305 ;
        RECT 46.805 -35.510 48.470 -35.340 ;
        RECT 46.250 -36.465 46.490 -36.115 ;
        RECT 47.470 -36.305 48.470 -35.510 ;
        RECT 46.320 -36.645 46.490 -36.465 ;
        RECT 45.400 -37.575 46.515 -37.530 ;
        RECT 43.985 -37.685 44.985 -37.575 ;
        RECT 43.100 -37.855 44.985 -37.685 ;
        RECT 45.400 -37.700 46.930 -37.575 ;
        RECT 42.530 -38.510 43.145 -38.340 ;
        RECT 42.975 -38.955 43.145 -38.510 ;
        RECT 43.985 -38.575 44.985 -37.855 ;
        RECT 45.930 -38.575 46.930 -37.700 ;
        RECT 42.560 -40.065 43.560 -39.650 ;
        RECT 42.045 -40.235 43.560 -40.065 ;
        RECT 42.560 -40.650 43.560 -40.235 ;
        RECT 40.160 -43.185 41.160 -42.185 ;
        RECT 83.315 -42.270 85.195 -42.100 ;
        RECT 85.735 -42.270 87.615 -42.100 ;
        RECT 6.470 -47.890 7.140 -47.720 ;
        RECT 7.680 -47.890 9.560 -47.720 ;
        RECT 10.100 -47.890 11.980 -47.720 ;
        RECT 7.605 -56.040 7.775 -51.480 ;
        RECT 8.280 -56.040 9.170 -55.725 ;
        RECT 7.605 -56.210 9.170 -56.040 ;
        RECT 7.605 -56.230 7.775 -56.210 ;
        RECT 8.280 -56.615 9.170 -56.210 ;
        RECT 17.495 -56.040 17.665 -51.480 ;
        RECT 18.180 -56.040 19.070 -55.725 ;
        RECT 17.495 -56.210 19.070 -56.040 ;
        RECT 17.495 -56.230 17.665 -56.210 ;
        RECT 18.180 -56.615 19.070 -56.210 ;
        RECT 27.330 -56.100 27.500 -51.525 ;
        RECT 27.860 -56.100 28.860 -55.540 ;
        RECT 36.890 -56.050 37.060 -51.480 ;
        RECT 37.485 -56.050 38.485 -55.945 ;
        RECT 27.330 -56.270 28.860 -56.100 ;
        RECT 36.870 -56.220 38.485 -56.050 ;
        RECT 36.890 -56.230 37.060 -56.220 ;
        RECT 27.330 -56.275 27.500 -56.270 ;
        RECT 27.860 -56.540 28.860 -56.270 ;
        RECT 5.315 -57.465 5.845 -56.935 ;
        RECT 15.280 -57.445 15.810 -56.915 ;
        RECT 37.485 -56.945 38.485 -56.220 ;
        RECT 43.415 -56.180 43.585 -47.190 ;
        RECT 45.975 -56.180 46.145 -47.190 ;
        RECT 48.535 -56.180 48.705 -47.190 ;
        RECT 51.095 -56.180 51.265 -47.190 ;
        RECT 53.655 -56.180 53.825 -47.190 ;
        RECT 61.060 -53.785 61.230 -47.170 ;
        RECT 61.060 -53.960 61.235 -53.785 ;
        RECT 63.620 -53.890 63.790 -47.170 ;
        RECT 66.180 -53.890 66.350 -47.170 ;
        RECT 68.740 -53.890 68.910 -47.170 ;
        RECT 71.300 -53.890 71.470 -47.170 ;
        RECT 63.620 -53.960 63.795 -53.890 ;
        RECT 66.180 -53.960 66.355 -53.890 ;
        RECT 68.740 -53.960 68.915 -53.890 ;
        RECT 71.300 -53.960 71.475 -53.890 ;
        RECT 54.235 -56.150 54.565 -56.075 ;
        RECT 55.400 -56.150 55.930 -55.995 ;
        RECT 54.235 -56.180 55.930 -56.150 ;
        RECT 43.415 -56.320 55.930 -56.180 ;
        RECT 59.110 -56.200 59.780 -55.590 ;
        RECT 43.415 -56.345 54.565 -56.320 ;
        RECT 43.415 -56.350 54.385 -56.345 ;
        RECT 43.415 -56.400 43.585 -56.350 ;
        RECT 55.400 -56.525 55.930 -56.320 ;
        RECT 61.065 -56.920 61.235 -53.960 ;
        RECT 25.040 -57.505 25.570 -56.975 ;
        RECT 34.740 -57.485 35.270 -56.955 ;
        RECT 60.635 -57.920 61.635 -56.920 ;
        RECT 63.625 -56.980 63.795 -53.960 ;
        RECT 66.185 -56.870 66.355 -53.960 ;
        RECT 68.745 -56.870 68.915 -53.960 ;
        RECT 71.305 -56.870 71.475 -53.960 ;
        RECT 63.205 -57.980 64.205 -56.980 ;
        RECT 65.710 -57.870 66.710 -56.870 ;
        RECT 68.320 -57.870 69.320 -56.870 ;
        RECT 70.805 -57.870 71.805 -56.870 ;
        RECT 74.635 -57.395 75.525 -57.110 ;
        RECT 76.265 -57.395 76.435 -51.210 ;
        RECT 74.635 -57.565 76.435 -57.395 ;
        RECT 74.635 -58.000 75.525 -57.565 ;
        RECT 76.265 -58.000 76.435 -57.565 ;
        RECT 77.175 -57.185 77.345 -51.210 ;
        RECT 78.065 -57.185 78.595 -57.005 ;
        RECT 77.175 -57.355 78.595 -57.185 ;
        RECT 77.175 -58.000 77.345 -57.355 ;
        RECT 78.065 -57.535 78.595 -57.355 ;
        RECT 2.475 -65.240 2.645 -65.055 ;
        RECT 3.280 -65.240 3.450 -60.760 ;
        RECT 2.475 -65.410 3.450 -65.240 ;
        RECT 2.475 -65.585 2.645 -65.410 ;
        RECT 3.280 -65.510 3.450 -65.410 ;
        RECT 7.560 -64.955 7.730 -60.760 ;
        RECT 8.260 -64.955 9.260 -64.585 ;
        RECT 7.560 -65.125 9.260 -64.955 ;
        RECT 7.560 -65.510 7.730 -65.125 ;
        RECT 8.260 -65.585 9.260 -65.125 ;
        RECT 12.415 -65.240 12.585 -65.055 ;
        RECT 13.155 -65.240 13.325 -60.760 ;
        RECT 12.415 -65.410 13.325 -65.240 ;
        RECT 12.415 -65.585 12.585 -65.410 ;
        RECT 13.155 -65.510 13.325 -65.410 ;
        RECT 17.435 -64.955 17.605 -60.760 ;
        RECT 18.155 -64.955 19.155 -64.585 ;
        RECT 17.435 -65.125 19.155 -64.955 ;
        RECT 17.435 -65.510 17.605 -65.125 ;
        RECT 18.155 -65.585 19.155 -65.125 ;
        RECT 22.080 -65.230 22.250 -65.055 ;
        RECT 23.095 -65.230 23.265 -60.760 ;
        RECT 22.080 -65.400 23.265 -65.230 ;
        RECT 22.080 -65.585 22.250 -65.400 ;
        RECT 23.095 -65.510 23.265 -65.400 ;
        RECT 27.375 -64.955 27.545 -60.760 ;
        RECT 28.010 -64.955 29.010 -64.585 ;
        RECT 27.375 -65.125 29.010 -64.955 ;
        RECT 27.375 -65.510 27.545 -65.125 ;
        RECT 28.010 -65.585 29.010 -65.125 ;
        RECT 31.595 -65.240 31.765 -65.055 ;
        RECT 32.515 -65.240 32.685 -60.760 ;
        RECT 31.595 -65.410 32.685 -65.240 ;
        RECT 31.595 -65.585 31.765 -65.410 ;
        RECT 32.515 -65.510 32.685 -65.410 ;
        RECT 36.795 -64.955 36.965 -60.760 ;
        RECT 37.185 -64.955 38.185 -64.585 ;
        RECT 36.795 -65.125 38.185 -64.955 ;
        RECT 36.795 -65.510 36.965 -65.125 ;
        RECT 37.185 -65.585 38.185 -65.125 ;
        RECT 7.105 -66.665 7.635 -66.135 ;
        RECT 13.300 -66.665 13.830 -66.135 ;
        RECT 23.305 -66.665 23.835 -66.135 ;
        RECT 32.570 -66.665 33.100 -66.135 ;
        RECT 43.525 -69.105 43.695 -59.545 ;
        RECT 45.345 -69.105 45.515 -59.545 ;
        RECT 47.165 -69.105 47.335 -59.545 ;
        RECT 48.985 -69.105 49.155 -59.545 ;
        RECT 50.805 -69.105 50.975 -59.545 ;
        RECT 52.625 -69.105 52.795 -59.545 ;
        RECT 53.550 -68.705 53.880 -68.435 ;
        RECT 53.635 -69.105 53.805 -68.705 ;
        RECT 54.445 -69.105 54.615 -59.545 ;
        RECT 59.320 -65.980 59.490 -59.290 ;
        RECT 59.305 -66.080 59.490 -65.980 ;
        RECT 59.305 -66.360 59.475 -66.080 ;
        RECT 59.305 -66.710 59.480 -66.360 ;
        RECT 59.310 -66.890 59.480 -66.710 ;
        RECT 60.230 -68.455 60.400 -59.290 ;
        RECT 61.140 -65.850 61.310 -59.290 ;
        RECT 61.125 -66.080 61.310 -65.850 ;
        RECT 61.125 -66.360 61.295 -66.080 ;
        RECT 61.125 -66.710 61.300 -66.360 ;
        RECT 61.130 -66.890 61.300 -66.710 ;
        RECT 62.050 -68.455 62.220 -59.290 ;
        RECT 62.960 -65.870 63.130 -59.290 ;
        RECT 62.945 -66.080 63.130 -65.870 ;
        RECT 62.945 -66.360 63.115 -66.080 ;
        RECT 62.945 -66.710 63.120 -66.360 ;
        RECT 62.950 -66.890 63.120 -66.710 ;
        RECT 63.870 -68.455 64.040 -59.290 ;
        RECT 64.780 -65.980 64.950 -59.290 ;
        RECT 64.780 -66.080 64.955 -65.980 ;
        RECT 64.785 -66.350 64.955 -66.080 ;
        RECT 64.770 -66.700 64.955 -66.350 ;
        RECT 64.770 -66.880 64.940 -66.700 ;
        RECT 65.690 -68.455 65.860 -59.290 ;
        RECT 66.600 -65.930 66.770 -59.290 ;
        RECT 66.600 -66.080 66.775 -65.930 ;
        RECT 66.605 -66.350 66.775 -66.080 ;
        RECT 66.590 -66.700 66.775 -66.350 ;
        RECT 66.590 -66.880 66.760 -66.700 ;
        RECT 67.510 -68.455 67.680 -59.290 ;
        RECT 68.420 -65.835 68.590 -59.290 ;
        RECT 68.405 -66.080 68.590 -65.835 ;
        RECT 68.405 -66.350 68.575 -66.080 ;
        RECT 68.405 -66.700 68.585 -66.350 ;
        RECT 68.415 -66.880 68.585 -66.700 ;
        RECT 69.330 -68.455 69.500 -59.290 ;
        RECT 70.240 -65.845 70.410 -59.290 ;
        RECT 70.225 -66.080 70.410 -65.845 ;
        RECT 70.225 -66.890 70.395 -66.080 ;
        RECT 71.150 -68.455 71.320 -59.290 ;
        RECT 72.060 -65.885 72.230 -59.290 ;
        RECT 72.045 -66.080 72.230 -65.885 ;
        RECT 72.045 -66.350 72.215 -66.080 ;
        RECT 72.045 -66.420 72.220 -66.350 ;
        RECT 71.930 -66.615 72.220 -66.420 ;
        RECT 72.050 -66.880 72.220 -66.615 ;
        RECT 55.345 -69.105 55.515 -68.890 ;
        RECT 43.525 -69.275 55.515 -69.105 ;
        RECT 55.345 -69.420 55.515 -69.275 ;
        RECT 59.750 -69.455 60.750 -68.455 ;
        RECT 61.635 -69.455 62.635 -68.455 ;
        RECT 63.460 -69.455 64.460 -68.455 ;
        RECT 65.335 -69.455 66.335 -68.455 ;
        RECT 67.155 -69.455 68.155 -68.455 ;
        RECT 68.895 -69.455 69.895 -68.455 ;
        RECT 70.730 -69.455 71.730 -68.455 ;
        RECT 58.755 -70.840 59.645 -69.950 ;
        RECT 2.475 -75.475 2.645 -75.290 ;
        RECT 3.280 -75.475 3.450 -70.910 ;
        RECT 2.475 -75.645 3.450 -75.475 ;
        RECT 2.475 -75.820 2.645 -75.645 ;
        RECT 3.280 -75.660 3.450 -75.645 ;
        RECT 7.560 -75.450 7.730 -70.910 ;
        RECT 8.200 -75.450 9.200 -75.080 ;
        RECT 7.560 -75.620 9.200 -75.450 ;
        RECT 7.560 -75.660 7.730 -75.620 ;
        RECT 8.200 -76.080 9.200 -75.620 ;
        RECT 12.435 -75.475 12.605 -75.290 ;
        RECT 13.175 -75.475 13.345 -70.910 ;
        RECT 12.435 -75.645 13.345 -75.475 ;
        RECT 12.435 -75.820 12.605 -75.645 ;
        RECT 13.175 -75.660 13.345 -75.645 ;
        RECT 17.455 -75.450 17.625 -70.910 ;
        RECT 18.110 -75.450 19.110 -75.080 ;
        RECT 17.455 -75.620 19.110 -75.450 ;
        RECT 17.455 -75.660 17.625 -75.620 ;
        RECT 18.110 -76.080 19.110 -75.620 ;
        RECT 22.205 -75.465 22.375 -75.290 ;
        RECT 23.220 -75.465 23.390 -70.910 ;
        RECT 22.205 -75.635 23.390 -75.465 ;
        RECT 22.205 -75.820 22.375 -75.635 ;
        RECT 23.220 -75.660 23.390 -75.635 ;
        RECT 27.500 -75.450 27.670 -70.910 ;
        RECT 28.125 -75.450 29.125 -75.080 ;
        RECT 27.500 -75.620 29.125 -75.450 ;
        RECT 27.500 -75.660 27.670 -75.620 ;
        RECT 28.125 -76.080 29.125 -75.620 ;
        RECT 31.640 -75.475 31.810 -75.290 ;
        RECT 32.420 -75.475 32.590 -70.910 ;
        RECT 31.640 -75.645 32.590 -75.475 ;
        RECT 31.640 -75.820 31.810 -75.645 ;
        RECT 32.420 -75.660 32.590 -75.645 ;
        RECT 36.700 -75.450 36.870 -70.910 ;
        RECT 74.940 -71.225 75.940 -70.895 ;
        RECT 76.440 -71.225 76.610 -64.660 ;
        RECT 74.940 -71.395 76.610 -71.225 ;
        RECT 74.940 -71.895 75.940 -71.395 ;
        RECT 76.440 -71.450 76.610 -71.395 ;
        RECT 77.350 -71.265 77.520 -64.660 ;
        RECT 84.525 -67.335 86.405 -67.165 ;
        RECT 86.945 -67.335 88.825 -67.165 ;
        RECT 77.985 -71.265 78.985 -70.895 ;
        RECT 77.350 -71.435 78.985 -71.265 ;
        RECT 77.350 -71.450 77.520 -71.435 ;
        RECT 77.985 -71.895 78.985 -71.435 ;
        RECT 42.750 -72.590 43.280 -72.060 ;
        RECT 48.085 -72.570 48.615 -72.040 ;
        RECT 56.570 -72.590 57.100 -72.060 ;
        RECT 62.140 -72.570 62.670 -72.040 ;
        RECT 37.330 -75.450 38.330 -75.080 ;
        RECT 36.700 -75.620 38.330 -75.450 ;
        RECT 36.700 -75.660 36.870 -75.620 ;
        RECT 37.330 -76.080 38.330 -75.620 ;
        RECT 7.075 -76.825 7.605 -76.295 ;
        RECT 17.005 -76.825 17.535 -76.295 ;
        RECT 27.055 -76.825 27.585 -76.295 ;
        RECT 32.475 -76.825 33.005 -76.295 ;
        RECT 5.110 -79.265 5.640 -78.735 ;
        RECT 15.220 -79.245 15.750 -78.715 ;
        RECT 25.295 -79.265 25.825 -78.735 ;
        RECT 34.495 -79.245 35.025 -78.715 ;
        RECT 43.870 -78.840 44.040 -73.230 ;
        RECT 44.505 -78.840 45.505 -78.470 ;
        RECT 43.870 -79.000 45.505 -78.840 ;
        RECT 50.560 -78.840 50.730 -73.230 ;
        RECT 51.195 -78.840 52.195 -78.470 ;
        RECT 57.250 -78.840 57.420 -73.230 ;
        RECT 57.860 -78.840 58.860 -78.470 ;
        RECT 63.890 -78.840 64.060 -73.230 ;
        RECT 68.715 -75.810 69.245 -75.280 ;
        RECT 75.050 -75.790 75.580 -75.260 ;
        RECT 81.075 -75.790 81.605 -75.260 ;
        RECT 87.420 -75.790 87.950 -75.260 ;
        RECT 64.485 -78.840 65.485 -78.470 ;
        RECT 50.560 -79.000 52.195 -78.840 ;
        RECT 43.890 -79.010 45.505 -79.000 ;
        RECT 50.580 -79.010 52.195 -79.000 ;
        RECT 57.245 -79.010 58.860 -78.840 ;
        RECT 63.870 -79.010 65.485 -78.840 ;
        RECT 44.505 -79.470 45.505 -79.010 ;
        RECT 51.195 -79.470 52.195 -79.010 ;
        RECT 57.860 -79.470 58.860 -79.010 ;
        RECT 64.485 -79.470 65.485 -79.010 ;
        RECT 7.615 -84.435 7.785 -79.925 ;
        RECT 8.235 -84.435 9.235 -84.065 ;
        RECT 7.615 -84.605 9.235 -84.435 ;
        RECT 7.615 -84.675 7.785 -84.605 ;
        RECT 8.235 -85.065 9.235 -84.605 ;
        RECT 17.430 -84.435 17.600 -79.925 ;
        RECT 18.145 -84.435 19.145 -84.065 ;
        RECT 17.430 -84.605 19.145 -84.435 ;
        RECT 17.430 -84.675 17.600 -84.605 ;
        RECT 18.145 -85.065 19.145 -84.605 ;
        RECT 27.590 -84.435 27.760 -79.925 ;
        RECT 28.300 -84.435 29.300 -84.065 ;
        RECT 27.590 -84.605 29.300 -84.435 ;
        RECT 27.590 -84.675 27.760 -84.605 ;
        RECT 28.300 -85.065 29.300 -84.605 ;
        RECT 36.655 -84.435 36.825 -79.925 ;
        RECT 70.090 -82.105 70.260 -76.525 ;
        RECT 70.705 -82.105 71.705 -81.735 ;
        RECT 70.090 -82.275 71.705 -82.105 ;
        RECT 70.090 -82.295 70.260 -82.275 ;
        RECT 70.705 -82.735 71.705 -82.275 ;
        RECT 76.785 -82.120 76.955 -76.525 ;
        RECT 77.410 -82.120 78.410 -81.750 ;
        RECT 82.900 -82.085 83.070 -76.525 ;
        RECT 83.505 -82.085 84.505 -81.715 ;
        RECT 76.785 -82.290 78.410 -82.120 ;
        RECT 82.890 -82.255 84.505 -82.085 ;
        RECT 89.305 -82.130 89.475 -76.525 ;
        RECT 89.910 -82.130 90.910 -81.760 ;
        RECT 76.785 -82.295 76.955 -82.290 ;
        RECT 77.410 -82.750 78.410 -82.290 ;
        RECT 82.900 -82.295 83.070 -82.255 ;
        RECT 83.505 -82.715 84.505 -82.255 ;
        RECT 89.295 -82.300 90.910 -82.130 ;
        RECT 89.910 -82.760 90.910 -82.300 ;
        RECT 37.305 -84.435 38.305 -84.065 ;
        RECT 36.655 -84.605 38.305 -84.435 ;
        RECT 36.655 -84.675 36.825 -84.605 ;
        RECT 37.305 -85.065 38.305 -84.605 ;
        RECT 68.300 -85.870 68.830 -85.340 ;
        RECT 75.005 -85.900 75.535 -85.370 ;
        RECT 81.095 -85.900 81.625 -85.370 ;
        RECT 87.570 -85.900 88.100 -85.370 ;
        RECT 70.090 -90.915 70.260 -86.650 ;
        RECT 70.715 -90.915 71.715 -90.545 ;
        RECT 70.090 -91.085 71.715 -90.915 ;
        RECT 70.090 -92.420 70.260 -91.085 ;
        RECT 70.715 -91.545 71.715 -91.085 ;
        RECT 76.785 -91.265 76.955 -86.650 ;
        RECT 77.420 -91.265 78.420 -90.895 ;
        RECT 76.785 -91.435 78.420 -91.265 ;
        RECT 76.785 -92.420 76.955 -91.435 ;
        RECT 77.420 -91.895 78.420 -91.435 ;
        RECT 82.900 -91.265 83.070 -86.650 ;
        RECT 83.535 -91.265 84.535 -90.895 ;
        RECT 82.900 -91.435 84.535 -91.265 ;
        RECT 82.900 -92.420 83.070 -91.435 ;
        RECT 83.535 -91.895 84.535 -91.435 ;
        RECT 89.305 -92.255 89.475 -86.650 ;
        RECT 89.930 -92.255 90.930 -91.885 ;
        RECT 89.305 -92.420 90.930 -92.255 ;
        RECT 89.315 -92.425 90.930 -92.420 ;
        RECT 89.930 -92.885 90.930 -92.425 ;
      LAYER met1 ;
        RECT 6.480 -7.085 8.340 -6.855 ;
        RECT 8.900 -7.085 10.760 -6.855 ;
        RECT 15.310 -13.660 15.950 -13.640 ;
        RECT 15.150 -14.560 16.110 -13.660 ;
        RECT 29.180 -14.530 30.180 -13.530 ;
        RECT 33.845 -13.630 34.485 -13.610 ;
        RECT 33.685 -14.530 34.645 -13.630 ;
        RECT 47.715 -14.500 48.715 -13.500 ;
        RECT 33.845 -14.550 34.485 -14.530 ;
        RECT 15.310 -14.580 15.950 -14.560 ;
        RECT 14.935 -16.065 15.935 -15.065 ;
        RECT 29.255 -15.230 29.895 -15.210 ;
        RECT 16.560 -15.590 17.200 -15.570 ;
        RECT 16.400 -16.490 17.360 -15.590 ;
        RECT 29.095 -16.130 30.055 -15.230 ;
        RECT 33.470 -16.035 34.470 -15.035 ;
        RECT 47.790 -15.200 48.430 -15.180 ;
        RECT 35.095 -15.560 35.735 -15.540 ;
        RECT 29.255 -16.150 29.895 -16.130 ;
        RECT 34.935 -16.460 35.895 -15.560 ;
        RECT 47.630 -16.100 48.590 -15.200 ;
        RECT 47.790 -16.120 48.430 -16.100 ;
        RECT 35.095 -16.480 35.735 -16.460 ;
        RECT 16.560 -16.510 17.200 -16.490 ;
        RECT 36.765 -16.610 37.405 -16.590 ;
        RECT 18.230 -16.640 18.870 -16.620 ;
        RECT 16.660 -17.970 17.660 -16.970 ;
        RECT 18.070 -17.540 19.030 -16.640 ;
        RECT 27.795 -17.310 28.435 -17.290 ;
        RECT 25.970 -17.515 26.610 -17.495 ;
        RECT 18.230 -17.560 18.870 -17.540 ;
        RECT 14.685 -18.205 15.335 -18.005 ;
        RECT 13.550 -18.345 15.335 -18.205 ;
        RECT 13.550 -37.375 13.690 -18.345 ;
        RECT 14.685 -18.595 15.335 -18.345 ;
        RECT 18.225 -19.000 19.225 -18.000 ;
        RECT 25.810 -18.415 26.770 -17.515 ;
        RECT 27.635 -18.210 28.595 -17.310 ;
        RECT 29.180 -17.685 30.180 -16.685 ;
        RECT 35.195 -17.940 36.195 -16.940 ;
        RECT 36.605 -17.510 37.565 -16.610 ;
        RECT 46.330 -17.280 46.970 -17.260 ;
        RECT 44.505 -17.485 45.145 -17.465 ;
        RECT 36.765 -17.530 37.405 -17.510 ;
        RECT 27.795 -18.230 28.435 -18.210 ;
        RECT 25.970 -18.435 26.610 -18.415 ;
        RECT 19.810 -18.755 20.450 -18.735 ;
        RECT 19.650 -19.655 20.610 -18.755 ;
        RECT 34.040 -18.925 34.690 -18.700 ;
        RECT 24.450 -19.620 25.090 -19.600 ;
        RECT 19.810 -19.675 20.450 -19.655 ;
        RECT 19.730 -21.350 20.730 -20.350 ;
        RECT 24.290 -20.520 25.250 -19.620 ;
        RECT 25.695 -19.955 26.695 -18.955 ;
        RECT 27.640 -19.955 28.640 -18.955 ;
        RECT 32.390 -19.065 34.690 -18.925 ;
        RECT 36.760 -18.970 37.760 -17.970 ;
        RECT 44.345 -18.385 45.305 -17.485 ;
        RECT 46.170 -18.180 47.130 -17.280 ;
        RECT 47.715 -17.655 48.715 -16.655 ;
        RECT 69.300 -17.750 69.950 -17.525 ;
        RECT 70.780 -17.750 71.420 -17.610 ;
        RECT 69.300 -17.890 71.420 -17.750 ;
        RECT 69.300 -18.115 69.950 -17.890 ;
        RECT 46.330 -18.200 46.970 -18.180 ;
        RECT 70.780 -18.190 71.420 -17.890 ;
        RECT 44.505 -18.405 45.145 -18.385 ;
        RECT 38.345 -18.725 38.985 -18.705 ;
        RECT 24.450 -20.540 25.090 -20.520 ;
        RECT 20.625 -21.955 21.265 -21.935 ;
        RECT 22.985 -21.955 23.625 -21.935 ;
        RECT 20.465 -22.855 21.425 -21.955 ;
        RECT 22.825 -22.855 23.785 -21.955 ;
        RECT 24.270 -22.030 25.270 -21.030 ;
        RECT 20.625 -22.875 21.265 -22.855 ;
        RECT 22.985 -22.875 23.625 -22.855 ;
        RECT 21.870 -24.565 22.870 -23.565 ;
        RECT 15.310 -31.990 15.950 -31.970 ;
        RECT 15.150 -32.890 16.110 -31.990 ;
        RECT 29.180 -32.860 30.180 -31.860 ;
        RECT 15.310 -32.910 15.950 -32.890 ;
        RECT 14.935 -34.395 15.935 -33.395 ;
        RECT 29.255 -33.560 29.895 -33.540 ;
        RECT 16.560 -33.920 17.200 -33.900 ;
        RECT 16.400 -34.820 17.360 -33.920 ;
        RECT 29.095 -34.460 30.055 -33.560 ;
        RECT 29.255 -34.480 29.895 -34.460 ;
        RECT 16.560 -34.840 17.200 -34.820 ;
        RECT 18.230 -34.970 18.870 -34.950 ;
        RECT 16.660 -36.300 17.660 -35.300 ;
        RECT 18.070 -35.870 19.030 -34.970 ;
        RECT 27.795 -35.640 28.435 -35.620 ;
        RECT 25.970 -35.845 26.610 -35.825 ;
        RECT 18.230 -35.890 18.870 -35.870 ;
        RECT 15.280 -37.375 15.930 -37.040 ;
        RECT 18.225 -37.330 19.225 -36.330 ;
        RECT 25.810 -36.745 26.770 -35.845 ;
        RECT 27.635 -36.540 28.595 -35.640 ;
        RECT 29.180 -36.015 30.180 -35.015 ;
        RECT 27.795 -36.560 28.435 -36.540 ;
        RECT 25.970 -36.765 26.610 -36.745 ;
        RECT 19.810 -37.085 20.450 -37.065 ;
        RECT 13.550 -37.515 15.930 -37.375 ;
        RECT 15.280 -37.630 15.930 -37.515 ;
        RECT 15.550 -44.655 15.690 -37.630 ;
        RECT 19.650 -37.985 20.610 -37.085 ;
        RECT 24.450 -37.950 25.090 -37.930 ;
        RECT 19.810 -38.005 20.450 -37.985 ;
        RECT 19.730 -39.680 20.730 -38.680 ;
        RECT 24.290 -38.850 25.250 -37.950 ;
        RECT 25.695 -38.285 26.695 -37.285 ;
        RECT 27.640 -38.285 28.640 -37.285 ;
        RECT 32.390 -37.625 32.530 -19.065 ;
        RECT 34.040 -19.290 34.690 -19.065 ;
        RECT 38.185 -19.625 39.145 -18.725 ;
        RECT 42.985 -19.590 43.625 -19.570 ;
        RECT 38.345 -19.645 38.985 -19.625 ;
        RECT 38.265 -21.320 39.265 -20.320 ;
        RECT 42.825 -20.490 43.785 -19.590 ;
        RECT 44.230 -19.925 45.230 -18.925 ;
        RECT 46.175 -19.925 47.175 -18.925 ;
        RECT 42.985 -20.510 43.625 -20.490 ;
        RECT 39.160 -21.925 39.800 -21.905 ;
        RECT 41.520 -21.925 42.160 -21.905 ;
        RECT 39.000 -22.825 39.960 -21.925 ;
        RECT 41.360 -22.825 42.320 -21.925 ;
        RECT 42.805 -22.000 43.805 -21.000 ;
        RECT 39.160 -22.845 39.800 -22.825 ;
        RECT 41.520 -22.845 42.160 -22.825 ;
        RECT 40.390 -24.535 41.390 -23.535 ;
        RECT 33.600 -32.280 34.240 -32.260 ;
        RECT 33.440 -33.180 34.400 -32.280 ;
        RECT 47.470 -33.150 48.470 -32.150 ;
        RECT 33.600 -33.200 34.240 -33.180 ;
        RECT 33.225 -34.635 34.225 -33.635 ;
        RECT 47.545 -33.850 48.185 -33.830 ;
        RECT 34.850 -34.210 35.490 -34.190 ;
        RECT 34.690 -35.110 35.650 -34.210 ;
        RECT 47.385 -34.750 48.345 -33.850 ;
        RECT 47.545 -34.770 48.185 -34.750 ;
        RECT 34.850 -35.130 35.490 -35.110 ;
        RECT 36.520 -35.260 37.160 -35.240 ;
        RECT 34.950 -36.590 35.950 -35.590 ;
        RECT 36.360 -36.160 37.320 -35.260 ;
        RECT 46.085 -35.930 46.725 -35.910 ;
        RECT 44.260 -36.135 44.900 -36.115 ;
        RECT 36.520 -36.180 37.160 -36.160 ;
        RECT 33.665 -37.625 34.315 -37.350 ;
        RECT 36.515 -37.620 37.515 -36.620 ;
        RECT 44.100 -37.035 45.060 -36.135 ;
        RECT 45.925 -36.830 46.885 -35.930 ;
        RECT 47.470 -36.305 48.470 -35.305 ;
        RECT 46.085 -36.850 46.725 -36.830 ;
        RECT 44.260 -37.055 44.900 -37.035 ;
        RECT 38.100 -37.375 38.740 -37.355 ;
        RECT 32.390 -37.765 34.435 -37.625 ;
        RECT 33.665 -37.940 34.435 -37.765 ;
        RECT 24.450 -38.870 25.090 -38.850 ;
        RECT 20.625 -40.285 21.265 -40.265 ;
        RECT 22.985 -40.285 23.625 -40.265 ;
        RECT 20.465 -41.185 21.425 -40.285 ;
        RECT 22.825 -41.185 23.785 -40.285 ;
        RECT 24.270 -40.360 25.270 -39.360 ;
        RECT 20.625 -41.205 21.265 -41.185 ;
        RECT 22.985 -41.205 23.625 -41.185 ;
        RECT 21.890 -42.895 22.890 -41.895 ;
        RECT 34.295 -44.655 34.435 -37.940 ;
        RECT 37.940 -38.275 38.900 -37.375 ;
        RECT 42.740 -38.240 43.380 -38.220 ;
        RECT 38.100 -38.295 38.740 -38.275 ;
        RECT 38.020 -39.970 39.020 -38.970 ;
        RECT 42.580 -39.140 43.540 -38.240 ;
        RECT 43.985 -38.575 44.985 -37.575 ;
        RECT 45.930 -38.575 46.930 -37.575 ;
        RECT 42.740 -39.160 43.380 -39.140 ;
        RECT 38.915 -40.575 39.555 -40.555 ;
        RECT 41.275 -40.575 41.915 -40.555 ;
        RECT 38.755 -41.475 39.715 -40.575 ;
        RECT 41.115 -41.475 42.075 -40.575 ;
        RECT 42.560 -40.650 43.560 -39.650 ;
        RECT 38.915 -41.495 39.555 -41.475 ;
        RECT 41.275 -41.495 41.915 -41.475 ;
        RECT 40.160 -43.185 41.160 -42.185 ;
        RECT 83.325 -42.300 85.185 -42.070 ;
        RECT 85.745 -42.300 87.605 -42.070 ;
        RECT 15.550 -44.795 56.205 -44.655 ;
        RECT 6.480 -47.725 7.130 -47.690 ;
        RECT 5.535 -47.865 7.130 -47.725 ;
        RECT 5.535 -48.095 5.675 -47.865 ;
        RECT 6.480 -47.920 7.130 -47.865 ;
        RECT 7.690 -47.920 9.550 -47.690 ;
        RECT 10.110 -47.920 11.970 -47.690 ;
        RECT 5.340 -48.675 5.980 -48.095 ;
        RECT 56.065 -54.955 56.205 -44.795 ;
        RECT 56.065 -55.095 56.685 -54.955 ;
        RECT 8.220 -56.645 9.230 -55.695 ;
        RECT 18.120 -56.645 19.130 -55.695 ;
        RECT 27.860 -56.540 28.860 -55.540 ;
        RECT 1.625 -57.115 2.265 -56.785 ;
        RECT 5.255 -57.115 5.905 -56.905 ;
        RECT 8.590 -57.115 8.730 -56.645 ;
        RECT 15.220 -57.115 15.870 -56.885 ;
        RECT 18.600 -57.115 18.740 -56.645 ;
        RECT 24.980 -57.115 25.630 -56.945 ;
        RECT 34.680 -57.115 35.330 -56.925 ;
        RECT 37.485 -56.945 38.485 -55.945 ;
        RECT 55.340 -56.555 55.990 -55.965 ;
        RECT 1.625 -57.255 35.330 -57.115 ;
        RECT 55.595 -57.230 55.735 -56.555 ;
        RECT 1.625 -57.365 2.265 -57.255 ;
        RECT 5.255 -57.495 5.905 -57.255 ;
        RECT 2.240 -64.870 2.880 -64.850 ;
        RECT 2.080 -65.770 3.040 -64.870 ;
        RECT 8.260 -65.585 9.260 -64.585 ;
        RECT 2.240 -65.790 2.880 -65.770 ;
        RECT 7.045 -66.335 7.695 -66.105 ;
        RECT 11.375 -66.335 11.515 -57.255 ;
        RECT 15.220 -57.475 15.870 -57.255 ;
        RECT 24.980 -57.535 25.630 -57.255 ;
        RECT 26.885 -57.270 27.025 -57.255 ;
        RECT 34.680 -57.515 35.330 -57.255 ;
        RECT 55.330 -57.810 55.970 -57.230 ;
        RECT 12.180 -64.870 12.820 -64.850 ;
        RECT 12.020 -65.770 12.980 -64.870 ;
        RECT 18.155 -65.585 19.155 -64.585 ;
        RECT 21.845 -64.870 22.485 -64.850 ;
        RECT 21.685 -65.770 22.645 -64.870 ;
        RECT 28.010 -65.585 29.010 -64.585 ;
        RECT 31.360 -64.870 32.000 -64.850 ;
        RECT 31.200 -65.770 32.160 -64.870 ;
        RECT 37.185 -65.585 38.185 -64.585 ;
        RECT 12.180 -65.790 12.820 -65.770 ;
        RECT 21.845 -65.790 22.485 -65.770 ;
        RECT 31.360 -65.790 32.000 -65.770 ;
        RECT 13.240 -66.335 13.890 -66.105 ;
        RECT 23.245 -66.330 23.895 -66.105 ;
        RECT 32.510 -66.330 33.160 -66.105 ;
        RECT 23.245 -66.335 33.160 -66.330 ;
        RECT 7.045 -66.470 33.160 -66.335 ;
        RECT 7.045 -66.475 23.895 -66.470 ;
        RECT 7.045 -66.695 7.695 -66.475 ;
        RECT 13.240 -66.695 13.890 -66.475 ;
        RECT 23.245 -66.695 23.895 -66.475 ;
        RECT 2.240 -75.105 2.880 -75.085 ;
        RECT 2.080 -76.005 3.040 -75.105 ;
        RECT 2.240 -76.025 2.880 -76.005 ;
        RECT 8.200 -76.080 9.200 -75.080 ;
        RECT 12.200 -75.105 12.840 -75.085 ;
        RECT 12.040 -76.005 13.000 -75.105 ;
        RECT 12.200 -76.025 12.840 -76.005 ;
        RECT 18.110 -76.080 19.110 -75.080 ;
        RECT 21.970 -75.105 22.610 -75.085 ;
        RECT 21.810 -76.005 22.770 -75.105 ;
        RECT 21.970 -76.025 22.610 -76.005 ;
        RECT 28.125 -76.080 29.125 -75.080 ;
        RECT 7.015 -76.490 7.665 -76.265 ;
        RECT 16.945 -76.490 17.595 -76.265 ;
        RECT 26.995 -76.490 27.645 -76.265 ;
        RECT 7.015 -76.500 27.645 -76.490 ;
        RECT 30.585 -76.500 30.725 -66.470 ;
        RECT 32.510 -66.695 33.160 -66.470 ;
        RECT 55.110 -68.705 55.750 -68.685 ;
        RECT 54.950 -69.605 55.910 -68.705 ;
        RECT 55.110 -69.625 55.750 -69.605 ;
        RECT 56.545 -70.380 56.685 -55.095 ;
        RECT 59.120 -56.190 59.770 -55.600 ;
        RECT 74.050 -56.180 74.690 -55.965 ;
        RECT 59.375 -57.230 59.515 -56.190 ;
        RECT 72.840 -56.480 74.690 -56.180 ;
        RECT 59.080 -57.810 59.720 -57.230 ;
        RECT 60.635 -57.920 61.635 -56.920 ;
        RECT 63.205 -57.980 64.205 -56.980 ;
        RECT 65.710 -57.870 66.710 -56.870 ;
        RECT 68.320 -57.870 69.320 -56.870 ;
        RECT 70.805 -57.870 71.805 -56.870 ;
        RECT 72.840 -57.195 73.140 -56.480 ;
        RECT 74.050 -56.545 74.690 -56.480 ;
        RECT 72.670 -57.775 73.310 -57.195 ;
        RECT 72.840 -60.505 73.140 -57.775 ;
        RECT 74.575 -58.030 75.585 -57.080 ;
        RECT 78.005 -57.565 78.655 -56.975 ;
        RECT 78.190 -60.505 78.490 -57.565 ;
        RECT 72.840 -60.805 78.490 -60.505 ;
        RECT 59.075 -66.175 59.715 -66.155 ;
        RECT 60.895 -66.175 61.535 -66.155 ;
        RECT 62.715 -66.175 63.355 -66.155 ;
        RECT 64.535 -66.165 65.175 -66.145 ;
        RECT 66.355 -66.165 66.995 -66.145 ;
        RECT 68.180 -66.165 68.820 -66.145 ;
        RECT 58.915 -67.075 59.875 -66.175 ;
        RECT 60.735 -67.075 61.695 -66.175 ;
        RECT 62.555 -67.075 63.515 -66.175 ;
        RECT 64.375 -67.065 65.335 -66.165 ;
        RECT 66.195 -67.065 67.155 -66.165 ;
        RECT 68.020 -67.065 68.980 -66.165 ;
        RECT 69.990 -66.175 70.630 -66.155 ;
        RECT 71.815 -66.165 72.455 -66.145 ;
        RECT 59.075 -67.095 59.715 -67.075 ;
        RECT 60.895 -67.095 61.535 -67.075 ;
        RECT 62.715 -67.095 63.355 -67.075 ;
        RECT 64.535 -67.085 65.175 -67.065 ;
        RECT 66.355 -67.085 66.995 -67.065 ;
        RECT 68.180 -67.085 68.820 -67.065 ;
        RECT 69.830 -67.075 70.790 -66.175 ;
        RECT 71.655 -67.065 72.615 -66.165 ;
        RECT 69.990 -67.095 70.630 -67.075 ;
        RECT 71.815 -67.085 72.455 -67.065 ;
        RECT 84.535 -67.365 86.395 -67.135 ;
        RECT 86.955 -67.365 88.815 -67.135 ;
        RECT 59.750 -69.455 60.750 -68.455 ;
        RECT 61.635 -69.455 62.635 -68.455 ;
        RECT 63.460 -69.455 64.460 -68.455 ;
        RECT 65.335 -69.455 66.335 -68.455 ;
        RECT 67.155 -69.455 68.155 -68.455 ;
        RECT 68.895 -69.455 69.895 -68.455 ;
        RECT 70.730 -69.455 71.730 -68.455 ;
        RECT 58.695 -70.325 59.705 -69.920 ;
        RECT 61.255 -70.325 61.895 -70.180 ;
        RECT 58.695 -70.380 61.895 -70.325 ;
        RECT 56.545 -70.465 61.895 -70.380 ;
        RECT 56.545 -70.520 59.705 -70.465 ;
        RECT 58.695 -70.870 59.705 -70.520 ;
        RECT 61.255 -70.760 61.895 -70.465 ;
        RECT 74.940 -71.895 75.940 -70.895 ;
        RECT 77.985 -71.895 78.985 -70.895 ;
        RECT 41.345 -72.255 41.985 -72.000 ;
        RECT 42.690 -72.240 43.340 -72.030 ;
        RECT 48.025 -72.240 48.675 -72.010 ;
        RECT 42.690 -72.255 48.675 -72.240 ;
        RECT 56.510 -72.240 57.160 -72.030 ;
        RECT 62.080 -72.240 62.730 -72.010 ;
        RECT 56.510 -72.255 62.730 -72.240 ;
        RECT 41.345 -72.380 62.730 -72.255 ;
        RECT 41.345 -72.395 43.340 -72.380 ;
        RECT 41.345 -72.580 41.985 -72.395 ;
        RECT 42.690 -72.620 43.340 -72.395 ;
        RECT 48.025 -72.395 57.160 -72.380 ;
        RECT 48.025 -72.600 48.675 -72.395 ;
        RECT 56.510 -72.620 57.160 -72.395 ;
        RECT 62.080 -72.600 62.730 -72.380 ;
        RECT 31.405 -75.105 32.045 -75.085 ;
        RECT 31.245 -76.005 32.205 -75.105 ;
        RECT 31.405 -76.025 32.045 -76.005 ;
        RECT 37.330 -76.080 38.330 -75.080 ;
        RECT 68.655 -75.460 69.305 -75.250 ;
        RECT 74.990 -75.455 75.640 -75.230 ;
        RECT 81.015 -75.455 81.665 -75.230 ;
        RECT 87.360 -75.455 88.010 -75.230 ;
        RECT 74.315 -75.460 92.535 -75.455 ;
        RECT 68.655 -75.595 92.535 -75.460 ;
        RECT 68.655 -75.600 74.460 -75.595 ;
        RECT 68.655 -75.840 69.305 -75.600 ;
        RECT 74.990 -75.820 75.640 -75.595 ;
        RECT 81.015 -75.820 81.665 -75.595 ;
        RECT 87.360 -75.820 88.010 -75.595 ;
        RECT 32.415 -76.500 33.065 -76.265 ;
        RECT 7.015 -76.630 33.065 -76.500 ;
        RECT 7.015 -76.855 7.665 -76.630 ;
        RECT 16.945 -76.855 17.595 -76.630 ;
        RECT 26.995 -76.640 33.065 -76.630 ;
        RECT 26.995 -76.855 27.645 -76.640 ;
        RECT 32.415 -76.855 33.065 -76.640 ;
        RECT 34.450 -78.500 35.090 -77.920 ;
        RECT 34.700 -78.685 34.840 -78.500 ;
        RECT 5.050 -78.915 5.700 -78.705 ;
        RECT 5.050 -78.930 14.125 -78.915 ;
        RECT 15.160 -78.930 15.810 -78.685 ;
        RECT 25.235 -78.930 25.885 -78.705 ;
        RECT 34.435 -78.930 35.085 -78.685 ;
        RECT 5.050 -79.055 35.085 -78.930 ;
        RECT 5.050 -79.295 5.700 -79.055 ;
        RECT 13.925 -79.070 35.085 -79.055 ;
        RECT 15.160 -79.275 15.810 -79.070 ;
        RECT 25.235 -79.295 25.885 -79.070 ;
        RECT 34.435 -79.275 35.085 -79.070 ;
        RECT 44.505 -79.470 45.505 -78.470 ;
        RECT 51.195 -79.470 52.195 -78.470 ;
        RECT 57.860 -79.470 58.860 -78.470 ;
        RECT 64.485 -79.470 65.485 -78.470 ;
        RECT 51.380 -83.020 52.020 -82.440 ;
        RECT 70.705 -82.735 71.705 -81.735 ;
        RECT 77.410 -82.750 78.410 -81.750 ;
        RECT 83.505 -82.715 84.505 -81.715 ;
        RECT 89.910 -82.760 90.910 -81.760 ;
        RECT 8.235 -85.065 9.235 -84.065 ;
        RECT 18.145 -85.065 19.145 -84.065 ;
        RECT 28.300 -85.065 29.300 -84.065 ;
        RECT 37.305 -85.065 38.305 -84.065 ;
        RECT 51.610 -85.570 51.750 -83.020 ;
        RECT 68.240 -85.570 68.890 -85.310 ;
        RECT 74.945 -85.565 75.595 -85.340 ;
        RECT 81.035 -85.565 81.685 -85.340 ;
        RECT 87.510 -85.565 88.160 -85.340 ;
        RECT 92.395 -85.565 92.535 -75.595 ;
        RECT 74.315 -85.570 92.535 -85.565 ;
        RECT 51.610 -85.705 92.535 -85.570 ;
        RECT 51.610 -85.710 74.460 -85.705 ;
        RECT 68.240 -85.900 68.890 -85.710 ;
        RECT 74.945 -85.930 75.595 -85.705 ;
        RECT 81.035 -85.930 81.685 -85.705 ;
        RECT 87.510 -85.930 88.160 -85.705 ;
        RECT 70.715 -91.545 71.715 -90.545 ;
        RECT 77.420 -91.895 78.420 -90.895 ;
        RECT 83.535 -91.895 84.535 -90.895 ;
        RECT 89.930 -92.885 90.930 -91.885 ;
      LAYER met2 ;
        RECT 15.150 -14.060 16.110 -13.660 ;
        RECT 14.250 -14.200 16.110 -14.060 ;
        RECT 14.250 -16.445 14.390 -14.200 ;
        RECT 15.150 -14.560 16.110 -14.200 ;
        RECT 29.095 -14.595 30.265 -13.465 ;
        RECT 33.685 -14.070 34.645 -13.630 ;
        RECT 32.785 -14.210 34.645 -14.070 ;
        RECT 14.850 -16.130 16.020 -15.000 ;
        RECT 16.400 -16.060 17.360 -15.590 ;
        RECT 29.095 -15.610 30.055 -15.230 ;
        RECT 29.095 -15.750 31.175 -15.610 ;
        RECT 16.400 -16.200 18.620 -16.060 ;
        RECT 29.095 -16.130 30.055 -15.750 ;
        RECT 16.400 -16.445 17.360 -16.200 ;
        RECT 14.250 -16.490 17.360 -16.445 ;
        RECT 14.250 -16.585 16.950 -16.490 ;
        RECT 14.250 -26.675 14.390 -16.585 ;
        RECT 18.480 -16.640 18.620 -16.200 ;
        RECT 16.575 -18.035 17.745 -16.905 ;
        RECT 18.070 -17.020 19.030 -16.640 ;
        RECT 18.070 -17.160 20.005 -17.020 ;
        RECT 18.070 -17.540 19.030 -17.160 ;
        RECT 18.140 -19.065 19.310 -17.935 ;
        RECT 19.865 -18.755 20.005 -17.160 ;
        RECT 25.810 -17.895 26.770 -17.515 ;
        RECT 24.735 -18.035 26.770 -17.895 ;
        RECT 19.650 -19.560 20.610 -18.755 ;
        RECT 18.825 -19.655 20.610 -19.560 ;
        RECT 24.735 -19.620 24.875 -18.035 ;
        RECT 25.810 -18.415 26.770 -18.035 ;
        RECT 27.635 -18.155 28.595 -17.310 ;
        RECT 29.095 -17.750 30.265 -16.620 ;
        RECT 27.635 -18.210 29.435 -18.155 ;
        RECT 28.045 -18.295 29.435 -18.210 ;
        RECT 18.825 -19.700 20.200 -19.655 ;
        RECT 18.825 -22.335 18.965 -19.700 ;
        RECT 24.290 -20.235 25.250 -19.620 ;
        RECT 25.610 -20.020 26.780 -18.890 ;
        RECT 27.555 -20.020 28.725 -18.890 ;
        RECT 29.295 -19.090 29.435 -18.295 ;
        RECT 31.035 -19.090 31.175 -15.750 ;
        RECT 29.295 -19.230 31.175 -19.090 ;
        RECT 32.785 -16.415 32.925 -14.210 ;
        RECT 33.685 -14.530 34.645 -14.210 ;
        RECT 47.630 -14.565 48.800 -13.435 ;
        RECT 33.385 -16.100 34.555 -14.970 ;
        RECT 34.935 -16.030 35.895 -15.560 ;
        RECT 47.630 -15.580 48.590 -15.200 ;
        RECT 47.630 -15.720 49.710 -15.580 ;
        RECT 34.935 -16.170 37.155 -16.030 ;
        RECT 47.630 -16.100 48.590 -15.720 ;
        RECT 34.935 -16.415 35.895 -16.170 ;
        RECT 32.785 -16.460 35.895 -16.415 ;
        RECT 32.785 -16.555 35.485 -16.460 ;
        RECT 19.645 -21.415 20.815 -20.285 ;
        RECT 24.290 -20.375 26.155 -20.235 ;
        RECT 24.290 -20.520 25.250 -20.375 ;
        RECT 26.015 -20.740 26.155 -20.375 ;
        RECT 29.295 -20.740 29.435 -19.230 ;
        RECT 26.015 -20.880 29.435 -20.740 ;
        RECT 20.465 -22.335 21.425 -21.955 ;
        RECT 22.825 -22.335 23.785 -21.955 ;
        RECT 24.185 -22.095 25.355 -20.965 ;
        RECT 18.825 -22.475 23.785 -22.335 ;
        RECT 20.465 -22.855 21.425 -22.475 ;
        RECT 22.825 -22.755 23.785 -22.475 ;
        RECT 26.015 -22.755 26.155 -20.880 ;
        RECT 22.825 -22.855 26.155 -22.755 ;
        RECT 23.235 -22.895 26.155 -22.855 ;
        RECT 21.785 -24.630 22.955 -23.500 ;
        RECT 32.785 -26.675 32.925 -16.555 ;
        RECT 37.015 -16.610 37.155 -16.170 ;
        RECT 35.110 -18.005 36.280 -16.875 ;
        RECT 36.605 -16.990 37.565 -16.610 ;
        RECT 36.605 -17.130 38.540 -16.990 ;
        RECT 36.605 -17.510 37.565 -17.130 ;
        RECT 36.675 -19.035 37.845 -17.905 ;
        RECT 38.400 -18.725 38.540 -17.130 ;
        RECT 44.345 -17.865 45.305 -17.485 ;
        RECT 43.270 -18.005 45.305 -17.865 ;
        RECT 38.185 -19.530 39.145 -18.725 ;
        RECT 37.360 -19.625 39.145 -19.530 ;
        RECT 43.270 -19.590 43.410 -18.005 ;
        RECT 44.345 -18.385 45.305 -18.005 ;
        RECT 46.170 -18.125 47.130 -17.280 ;
        RECT 47.630 -17.720 48.800 -16.590 ;
        RECT 46.170 -18.180 47.970 -18.125 ;
        RECT 46.580 -18.265 47.970 -18.180 ;
        RECT 37.360 -19.670 38.735 -19.625 ;
        RECT 37.360 -22.305 37.500 -19.670 ;
        RECT 42.825 -20.205 43.785 -19.590 ;
        RECT 44.145 -19.990 45.315 -18.860 ;
        RECT 46.090 -19.990 47.260 -18.860 ;
        RECT 47.830 -19.060 47.970 -18.265 ;
        RECT 49.570 -19.060 49.710 -15.720 ;
        RECT 70.780 -18.200 71.420 -17.600 ;
        RECT 47.830 -19.200 49.710 -19.060 ;
        RECT 38.180 -21.385 39.350 -20.255 ;
        RECT 42.825 -20.345 44.690 -20.205 ;
        RECT 42.825 -20.490 43.785 -20.345 ;
        RECT 44.550 -20.710 44.690 -20.345 ;
        RECT 47.830 -20.710 47.970 -19.200 ;
        RECT 44.550 -20.850 47.970 -20.710 ;
        RECT 39.000 -22.305 39.960 -21.925 ;
        RECT 41.360 -22.305 42.320 -21.925 ;
        RECT 42.720 -22.065 43.890 -20.935 ;
        RECT 37.360 -22.445 42.320 -22.305 ;
        RECT 39.000 -22.825 39.960 -22.445 ;
        RECT 41.360 -22.725 42.320 -22.445 ;
        RECT 44.550 -22.725 44.690 -20.850 ;
        RECT 41.360 -22.825 44.690 -22.725 ;
        RECT 41.770 -22.865 44.690 -22.825 ;
        RECT 40.305 -24.600 41.475 -23.470 ;
        RECT 14.250 -26.815 32.925 -26.675 ;
        RECT 14.250 -32.430 14.390 -26.815 ;
        RECT 15.150 -32.430 16.110 -31.990 ;
        RECT 14.250 -32.570 16.110 -32.430 ;
        RECT 14.250 -34.775 14.390 -32.570 ;
        RECT 15.150 -32.890 16.110 -32.570 ;
        RECT 29.095 -32.925 30.265 -31.795 ;
        RECT 32.785 -32.835 32.925 -26.815 ;
        RECT 71.030 -27.250 71.170 -18.200 ;
        RECT 50.990 -27.390 71.170 -27.250 ;
        RECT 33.440 -32.835 34.400 -32.280 ;
        RECT 32.785 -32.975 34.400 -32.835 ;
        RECT 14.850 -34.460 16.020 -33.330 ;
        RECT 16.400 -34.390 17.360 -33.920 ;
        RECT 29.095 -33.940 30.055 -33.560 ;
        RECT 29.095 -34.080 31.175 -33.940 ;
        RECT 16.400 -34.530 18.620 -34.390 ;
        RECT 29.095 -34.460 30.055 -34.080 ;
        RECT 16.400 -34.775 17.360 -34.530 ;
        RECT 14.250 -34.820 17.360 -34.775 ;
        RECT 14.250 -34.915 16.950 -34.820 ;
        RECT 18.480 -34.970 18.620 -34.530 ;
        RECT 16.575 -36.365 17.745 -35.235 ;
        RECT 18.070 -35.350 19.030 -34.970 ;
        RECT 18.070 -35.490 20.005 -35.350 ;
        RECT 18.070 -35.870 19.030 -35.490 ;
        RECT 18.140 -37.395 19.310 -36.265 ;
        RECT 19.865 -37.085 20.005 -35.490 ;
        RECT 25.810 -36.225 26.770 -35.845 ;
        RECT 24.735 -36.365 26.770 -36.225 ;
        RECT 19.650 -37.890 20.610 -37.085 ;
        RECT 18.825 -37.985 20.610 -37.890 ;
        RECT 24.735 -37.950 24.875 -36.365 ;
        RECT 25.810 -36.745 26.770 -36.365 ;
        RECT 27.635 -36.485 28.595 -35.640 ;
        RECT 29.095 -36.080 30.265 -34.950 ;
        RECT 27.635 -36.540 29.435 -36.485 ;
        RECT 28.045 -36.625 29.435 -36.540 ;
        RECT 18.825 -38.030 20.200 -37.985 ;
        RECT 18.825 -40.665 18.965 -38.030 ;
        RECT 24.290 -38.565 25.250 -37.950 ;
        RECT 25.610 -38.350 26.780 -37.220 ;
        RECT 27.555 -38.350 28.725 -37.220 ;
        RECT 29.295 -37.420 29.435 -36.625 ;
        RECT 31.035 -37.420 31.175 -34.080 ;
        RECT 32.785 -34.850 32.925 -32.975 ;
        RECT 33.440 -33.180 34.400 -32.975 ;
        RECT 47.385 -33.215 48.555 -32.085 ;
        RECT 33.140 -34.700 34.310 -33.570 ;
        RECT 34.690 -34.680 35.650 -34.210 ;
        RECT 47.385 -34.230 48.345 -33.850 ;
        RECT 50.990 -34.190 51.130 -27.390 ;
        RECT 49.935 -34.230 51.130 -34.190 ;
        RECT 47.385 -34.330 51.130 -34.230 ;
        RECT 47.385 -34.370 50.075 -34.330 ;
        RECT 34.690 -34.820 36.910 -34.680 ;
        RECT 47.385 -34.750 48.345 -34.370 ;
        RECT 34.690 -34.850 35.650 -34.820 ;
        RECT 32.785 -34.990 35.650 -34.850 ;
        RECT 34.690 -35.110 35.650 -34.990 ;
        RECT 36.770 -35.260 36.910 -34.820 ;
        RECT 34.865 -36.655 36.035 -35.525 ;
        RECT 36.360 -35.640 37.320 -35.260 ;
        RECT 36.360 -35.780 38.295 -35.640 ;
        RECT 36.360 -36.160 37.320 -35.780 ;
        RECT 29.295 -37.560 31.175 -37.420 ;
        RECT 19.645 -39.745 20.815 -38.615 ;
        RECT 24.290 -38.705 26.155 -38.565 ;
        RECT 24.290 -38.850 25.250 -38.705 ;
        RECT 26.015 -39.070 26.155 -38.705 ;
        RECT 29.295 -39.070 29.435 -37.560 ;
        RECT 36.430 -37.685 37.600 -36.555 ;
        RECT 38.155 -37.375 38.295 -35.780 ;
        RECT 44.100 -36.515 45.060 -36.135 ;
        RECT 43.400 -36.655 45.060 -36.515 ;
        RECT 37.940 -38.180 38.900 -37.375 ;
        RECT 26.015 -39.210 29.435 -39.070 ;
        RECT 37.115 -38.275 38.900 -38.180 ;
        RECT 43.400 -38.240 43.540 -36.655 ;
        RECT 44.100 -37.035 45.060 -36.655 ;
        RECT 45.925 -36.830 46.885 -35.930 ;
        RECT 47.385 -36.370 48.555 -35.240 ;
        RECT 46.335 -36.980 46.475 -36.830 ;
        RECT 46.335 -37.120 47.675 -36.980 ;
        RECT 37.115 -38.320 38.490 -38.275 ;
        RECT 20.465 -40.665 21.425 -40.285 ;
        RECT 22.825 -40.665 23.785 -40.285 ;
        RECT 24.185 -40.425 25.355 -39.295 ;
        RECT 18.825 -40.805 23.785 -40.665 ;
        RECT 20.465 -41.185 21.425 -40.805 ;
        RECT 22.825 -41.085 23.785 -40.805 ;
        RECT 26.015 -41.085 26.155 -39.210 ;
        RECT 22.825 -41.185 26.155 -41.085 ;
        RECT 37.115 -40.955 37.255 -38.320 ;
        RECT 42.580 -38.855 43.540 -38.240 ;
        RECT 43.900 -38.640 45.070 -37.510 ;
        RECT 45.845 -38.640 47.015 -37.510 ;
        RECT 47.535 -37.710 47.675 -37.120 ;
        RECT 49.700 -37.710 49.840 -34.370 ;
        RECT 47.535 -37.850 49.840 -37.710 ;
        RECT 37.935 -40.035 39.105 -38.905 ;
        RECT 42.580 -38.995 44.820 -38.855 ;
        RECT 42.580 -39.140 43.540 -38.995 ;
        RECT 44.680 -39.190 44.820 -38.995 ;
        RECT 47.535 -39.190 47.675 -37.850 ;
        RECT 44.680 -39.330 47.675 -39.190 ;
        RECT 38.755 -40.955 39.715 -40.575 ;
        RECT 41.115 -40.955 42.075 -40.575 ;
        RECT 42.475 -40.715 43.645 -39.585 ;
        RECT 37.115 -41.095 42.075 -40.955 ;
        RECT 23.235 -41.225 26.155 -41.185 ;
        RECT 38.755 -41.475 39.715 -41.095 ;
        RECT 41.115 -41.375 42.075 -41.095 ;
        RECT 44.680 -41.375 44.820 -39.330 ;
        RECT 41.115 -41.475 44.820 -41.375 ;
        RECT 41.525 -41.515 44.820 -41.475 ;
        RECT 21.805 -42.960 22.975 -41.830 ;
        RECT 40.075 -43.250 41.245 -42.120 ;
        RECT 44.680 -45.450 44.820 -41.515 ;
        RECT 44.680 -45.470 73.265 -45.450 ;
        RECT 44.680 -45.590 74.385 -45.470 ;
        RECT 73.125 -45.610 74.385 -45.590 ;
        RECT 1.225 -48.095 5.730 -48.025 ;
        RECT 1.225 -48.165 5.980 -48.095 ;
        RECT 1.225 -66.560 1.365 -48.165 ;
        RECT 5.340 -48.675 5.980 -48.165 ;
        RECT 27.775 -56.605 28.945 -55.475 ;
        RECT 1.560 -57.440 2.330 -56.710 ;
        RECT 37.400 -57.010 38.570 -55.880 ;
        RECT 74.245 -55.965 74.385 -45.610 ;
        RECT 74.050 -56.545 74.690 -55.965 ;
        RECT 55.265 -57.885 56.035 -57.155 ;
        RECT 59.015 -57.885 59.785 -57.155 ;
        RECT 60.550 -57.985 61.720 -56.855 ;
        RECT 63.120 -58.045 64.290 -56.915 ;
        RECT 65.625 -57.935 66.795 -56.805 ;
        RECT 68.235 -57.935 69.405 -56.805 ;
        RECT 70.720 -57.935 71.890 -56.805 ;
        RECT 72.605 -57.850 73.375 -57.120 ;
        RECT 74.495 -58.120 75.665 -56.990 ;
        RECT 2.080 -65.770 3.040 -64.870 ;
        RECT 8.175 -65.650 9.345 -64.520 ;
        RECT 12.020 -65.770 12.980 -64.870 ;
        RECT 18.070 -65.650 19.240 -64.520 ;
        RECT 21.685 -65.770 22.645 -64.870 ;
        RECT 27.925 -65.650 29.095 -64.520 ;
        RECT 31.200 -65.770 32.160 -64.870 ;
        RECT 37.100 -65.650 38.270 -64.520 ;
        RECT 2.490 -66.560 2.630 -65.770 ;
        RECT 12.520 -66.560 12.660 -65.770 ;
        RECT 22.095 -66.560 22.235 -65.770 ;
        RECT 31.655 -66.560 31.795 -65.770 ;
        RECT 1.225 -66.700 31.795 -66.560 ;
        RECT 58.915 -66.575 59.875 -66.175 ;
        RECT 1.225 -76.745 1.365 -66.700 ;
        RECT 57.420 -66.715 59.875 -66.575 ;
        RECT 54.950 -69.085 55.910 -68.705 ;
        RECT 57.420 -69.085 57.560 -66.715 ;
        RECT 58.915 -67.075 59.875 -66.715 ;
        RECT 60.735 -67.075 61.695 -66.175 ;
        RECT 62.555 -67.075 63.515 -66.175 ;
        RECT 64.375 -67.065 65.335 -66.165 ;
        RECT 66.195 -67.065 67.155 -66.165 ;
        RECT 68.020 -67.065 68.980 -66.165 ;
        RECT 59.315 -67.550 59.455 -67.075 ;
        RECT 61.295 -67.550 61.435 -67.075 ;
        RECT 62.945 -67.550 63.085 -67.075 ;
        RECT 64.810 -67.550 64.950 -67.065 ;
        RECT 66.615 -67.550 66.755 -67.065 ;
        RECT 68.440 -67.550 68.580 -67.065 ;
        RECT 69.830 -67.075 70.790 -66.175 ;
        RECT 71.655 -67.065 72.615 -66.165 ;
        RECT 70.245 -67.550 70.385 -67.075 ;
        RECT 72.065 -67.550 72.205 -67.065 ;
        RECT 59.315 -67.690 72.205 -67.550 ;
        RECT 54.950 -69.225 57.560 -69.085 ;
        RECT 54.950 -69.605 55.910 -69.225 ;
        RECT 59.665 -69.520 60.835 -68.390 ;
        RECT 61.550 -69.520 62.720 -68.390 ;
        RECT 63.375 -69.520 64.545 -68.390 ;
        RECT 65.250 -69.520 66.420 -68.390 ;
        RECT 67.070 -69.520 68.240 -68.390 ;
        RECT 68.810 -69.520 69.980 -68.390 ;
        RECT 70.645 -69.520 71.815 -68.390 ;
        RECT 60.990 -71.035 62.160 -69.905 ;
        RECT 41.280 -72.655 42.050 -71.925 ;
        RECT 74.855 -71.960 76.025 -70.830 ;
        RECT 77.900 -71.960 79.070 -70.830 ;
        RECT 2.080 -76.005 3.040 -75.105 ;
        RECT 2.490 -76.745 2.630 -76.005 ;
        RECT 8.115 -76.145 9.285 -75.015 ;
        RECT 12.040 -76.005 13.000 -75.105 ;
        RECT 12.540 -76.745 12.680 -76.005 ;
        RECT 18.025 -76.145 19.195 -75.015 ;
        RECT 21.810 -76.005 22.770 -75.105 ;
        RECT 22.220 -76.745 22.360 -76.005 ;
        RECT 28.040 -76.145 29.210 -75.015 ;
        RECT 31.245 -76.005 32.205 -75.105 ;
        RECT 31.685 -76.745 31.825 -76.005 ;
        RECT 37.245 -76.145 38.415 -75.015 ;
        RECT 1.225 -76.885 31.825 -76.745 ;
        RECT 12.540 -76.895 12.680 -76.885 ;
        RECT 22.220 -76.895 22.360 -76.885 ;
        RECT 34.385 -78.575 35.155 -77.845 ;
        RECT 44.420 -79.535 45.590 -78.405 ;
        RECT 51.110 -79.535 52.280 -78.405 ;
        RECT 57.775 -79.535 58.945 -78.405 ;
        RECT 64.400 -79.535 65.570 -78.405 ;
        RECT 51.315 -83.095 52.085 -82.365 ;
        RECT 70.620 -82.800 71.790 -81.670 ;
        RECT 77.325 -82.815 78.495 -81.685 ;
        RECT 83.420 -82.780 84.590 -81.650 ;
        RECT 89.825 -82.825 90.995 -81.695 ;
        RECT 8.150 -85.130 9.320 -84.000 ;
        RECT 18.060 -85.130 19.230 -84.000 ;
        RECT 28.215 -85.130 29.385 -84.000 ;
        RECT 37.220 -85.130 38.390 -84.000 ;
        RECT 70.630 -91.610 71.800 -90.480 ;
        RECT 77.335 -91.960 78.505 -90.830 ;
        RECT 83.450 -91.960 84.620 -90.830 ;
        RECT 89.845 -92.950 91.015 -91.820 ;
      LAYER met3 ;
        RECT 29.095 -13.680 30.265 -13.465 ;
        RECT 47.630 -13.640 48.800 -13.435 ;
        RECT 29.095 -14.380 31.270 -13.680 ;
        RECT 29.095 -14.595 30.265 -14.380 ;
        RECT 14.850 -16.130 16.020 -15.000 ;
        RECT 15.045 -17.120 15.745 -16.130 ;
        RECT 29.095 -16.705 30.265 -16.620 ;
        RECT 30.570 -16.705 31.270 -14.380 ;
        RECT 47.630 -14.340 49.905 -13.640 ;
        RECT 47.630 -14.565 48.800 -14.340 ;
        RECT 33.385 -16.100 34.555 -14.970 ;
        RECT 16.575 -17.120 17.745 -16.905 ;
        RECT 15.045 -17.820 17.745 -17.120 ;
        RECT 29.095 -17.405 31.270 -16.705 ;
        RECT 33.580 -17.090 34.280 -16.100 ;
        RECT 47.630 -16.805 48.800 -16.590 ;
        RECT 49.205 -16.805 49.905 -14.340 ;
        RECT 35.110 -17.090 36.280 -16.875 ;
        RECT 29.095 -17.750 30.265 -17.405 ;
        RECT 16.575 -18.035 17.745 -17.820 ;
        RECT 16.800 -18.370 17.500 -18.035 ;
        RECT 18.140 -18.150 19.310 -17.935 ;
        RECT 18.070 -18.370 19.310 -18.150 ;
        RECT 16.800 -19.065 19.310 -18.370 ;
        RECT 16.800 -19.070 18.770 -19.065 ;
        RECT 18.070 -20.500 18.770 -19.070 ;
        RECT 25.610 -19.105 26.780 -18.890 ;
        RECT 27.555 -19.105 28.725 -18.890 ;
        RECT 25.610 -19.240 28.725 -19.105 ;
        RECT 29.450 -19.240 30.150 -17.750 ;
        RECT 33.580 -17.790 36.280 -17.090 ;
        RECT 47.630 -17.505 49.905 -16.805 ;
        RECT 47.630 -17.720 48.800 -17.505 ;
        RECT 35.110 -18.005 36.280 -17.790 ;
        RECT 35.335 -18.345 36.035 -18.005 ;
        RECT 36.675 -18.335 37.845 -17.905 ;
        RECT 36.545 -18.345 37.845 -18.335 ;
        RECT 35.335 -19.035 37.845 -18.345 ;
        RECT 35.335 -19.045 37.260 -19.035 ;
        RECT 25.610 -19.805 30.150 -19.240 ;
        RECT 25.610 -20.020 26.895 -19.805 ;
        RECT 27.555 -19.940 30.150 -19.805 ;
        RECT 27.555 -20.020 28.725 -19.940 ;
        RECT 19.645 -20.500 20.815 -20.285 ;
        RECT 18.070 -21.200 20.815 -20.500 ;
        RECT 19.645 -21.415 20.815 -21.200 ;
        RECT 24.185 -21.040 25.355 -20.965 ;
        RECT 26.195 -21.040 26.895 -20.020 ;
        RECT 19.940 -23.670 20.640 -21.415 ;
        RECT 24.185 -21.740 26.895 -21.040 ;
        RECT 24.185 -22.095 25.355 -21.740 ;
        RECT 21.785 -23.655 22.955 -23.500 ;
        RECT 24.420 -23.655 25.120 -22.095 ;
        RECT 21.785 -23.670 25.120 -23.655 ;
        RECT 19.940 -24.355 25.120 -23.670 ;
        RECT 19.940 -24.370 22.955 -24.355 ;
        RECT 21.785 -24.630 22.955 -24.370 ;
        RECT 29.450 -26.895 30.150 -19.940 ;
        RECT 36.545 -20.685 37.245 -19.045 ;
        RECT 44.145 -19.075 45.315 -18.860 ;
        RECT 46.090 -19.075 47.260 -18.860 ;
        RECT 44.145 -19.210 47.260 -19.075 ;
        RECT 48.085 -19.210 48.785 -17.720 ;
        RECT 44.145 -19.775 48.785 -19.210 ;
        RECT 44.145 -19.990 45.430 -19.775 ;
        RECT 46.090 -19.910 48.785 -19.775 ;
        RECT 46.090 -19.990 47.260 -19.910 ;
        RECT 38.180 -20.685 39.350 -20.255 ;
        RECT 36.545 -21.385 39.350 -20.685 ;
        RECT 42.720 -21.010 43.890 -20.935 ;
        RECT 44.730 -21.010 45.430 -19.990 ;
        RECT 38.415 -23.855 39.115 -21.385 ;
        RECT 42.720 -21.710 45.430 -21.010 ;
        RECT 42.720 -22.065 43.890 -21.710 ;
        RECT 40.305 -23.855 41.475 -23.470 ;
        RECT 42.955 -23.855 43.655 -22.065 ;
        RECT 38.415 -24.555 43.655 -23.855 ;
        RECT 40.305 -24.600 41.475 -24.555 ;
        RECT 48.085 -26.895 48.785 -19.910 ;
        RECT 29.450 -27.595 48.785 -26.895 ;
        RECT 29.450 -31.795 30.150 -27.595 ;
        RECT 48.085 -27.785 48.785 -27.595 ;
        RECT 49.450 -27.785 50.230 -27.710 ;
        RECT 48.085 -28.430 50.230 -27.785 ;
        RECT 48.085 -28.485 50.190 -28.430 ;
        RECT 29.095 -32.000 30.265 -31.795 ;
        RECT 29.095 -32.700 31.290 -32.000 ;
        RECT 48.085 -32.085 48.785 -28.485 ;
        RECT 75.630 -28.940 98.080 -6.485 ;
        RECT 29.095 -32.925 30.265 -32.700 ;
        RECT 14.850 -34.460 16.020 -33.330 ;
        RECT 15.045 -35.450 15.745 -34.460 ;
        RECT 29.095 -35.165 30.265 -34.950 ;
        RECT 30.590 -35.165 31.290 -32.700 ;
        RECT 47.385 -32.290 48.785 -32.085 ;
        RECT 47.385 -33.000 49.670 -32.290 ;
        RECT 47.385 -33.215 48.555 -33.000 ;
        RECT 33.140 -34.700 34.310 -33.570 ;
        RECT 16.575 -35.450 17.745 -35.235 ;
        RECT 15.045 -36.150 17.745 -35.450 ;
        RECT 29.095 -35.865 31.290 -35.165 ;
        RECT 33.335 -35.740 34.035 -34.700 ;
        RECT 47.385 -35.455 48.555 -35.240 ;
        RECT 48.970 -35.455 49.670 -33.000 ;
        RECT 34.865 -35.740 36.035 -35.525 ;
        RECT 29.095 -36.080 30.265 -35.865 ;
        RECT 16.575 -36.365 17.745 -36.150 ;
        RECT 16.800 -36.785 17.500 -36.365 ;
        RECT 18.140 -36.785 19.310 -36.265 ;
        RECT 16.800 -37.395 19.310 -36.785 ;
        RECT 16.800 -37.485 18.855 -37.395 ;
        RECT 18.155 -38.830 18.855 -37.485 ;
        RECT 25.610 -37.435 26.780 -37.220 ;
        RECT 27.555 -37.435 28.725 -37.220 ;
        RECT 25.610 -37.570 28.725 -37.435 ;
        RECT 29.470 -37.570 30.170 -36.080 ;
        RECT 33.335 -36.440 36.035 -35.740 ;
        RECT 47.385 -36.155 49.670 -35.455 ;
        RECT 47.385 -36.370 48.555 -36.155 ;
        RECT 34.865 -36.655 36.035 -36.440 ;
        RECT 25.610 -38.135 30.170 -37.570 ;
        RECT 35.090 -36.970 35.790 -36.655 ;
        RECT 36.430 -36.965 37.600 -36.555 ;
        RECT 36.300 -36.970 37.600 -36.965 ;
        RECT 35.090 -37.670 37.600 -36.970 ;
        RECT 25.610 -38.350 27.035 -38.135 ;
        RECT 27.555 -38.270 30.170 -38.135 ;
        RECT 36.300 -37.685 37.600 -37.670 ;
        RECT 27.555 -38.350 28.725 -38.270 ;
        RECT 19.645 -38.830 20.815 -38.615 ;
        RECT 18.155 -39.530 20.815 -38.830 ;
        RECT 19.645 -39.745 20.815 -39.530 ;
        RECT 24.185 -39.370 25.355 -39.295 ;
        RECT 26.335 -39.370 27.035 -38.350 ;
        RECT 20.025 -42.000 20.725 -39.745 ;
        RECT 24.185 -40.070 27.035 -39.370 ;
        RECT 36.300 -39.315 37.000 -37.685 ;
        RECT 43.900 -37.725 45.070 -37.510 ;
        RECT 45.845 -37.725 47.015 -37.510 ;
        RECT 43.900 -37.860 47.015 -37.725 ;
        RECT 47.850 -37.860 48.550 -36.370 ;
        RECT 43.900 -38.425 48.550 -37.860 ;
        RECT 43.900 -38.640 45.415 -38.425 ;
        RECT 45.845 -38.560 48.550 -38.425 ;
        RECT 45.845 -38.640 47.015 -38.560 ;
        RECT 37.935 -39.315 39.105 -38.905 ;
        RECT 36.300 -40.015 39.105 -39.315 ;
        RECT 37.935 -40.035 39.105 -40.015 ;
        RECT 42.475 -39.660 43.645 -39.585 ;
        RECT 44.715 -39.660 45.415 -38.640 ;
        RECT 24.185 -40.425 25.355 -40.070 ;
        RECT 21.805 -41.985 22.975 -41.830 ;
        RECT 24.560 -41.985 25.260 -40.425 ;
        RECT 21.805 -42.000 25.260 -41.985 ;
        RECT 20.025 -42.685 25.260 -42.000 ;
        RECT 38.170 -42.485 38.870 -40.035 ;
        RECT 42.475 -40.360 45.415 -39.660 ;
        RECT 42.475 -40.715 43.645 -40.360 ;
        RECT 40.075 -42.485 41.245 -42.120 ;
        RECT 42.940 -42.485 43.640 -40.715 ;
        RECT 20.025 -42.700 22.975 -42.685 ;
        RECT 21.805 -42.960 22.975 -42.700 ;
        RECT 38.170 -43.185 43.640 -42.485 ;
        RECT 40.075 -43.250 41.245 -43.185 ;
        RECT 27.775 -56.605 28.945 -55.475 ;
        RECT 1.560 -57.440 2.330 -56.710 ;
        RECT 1.680 -86.500 1.980 -57.440 ;
        RECT 28.175 -57.855 28.475 -56.605 ;
        RECT 37.400 -57.010 38.570 -55.880 ;
        RECT 37.865 -57.855 38.165 -57.010 ;
        RECT 28.175 -58.155 39.015 -57.855 ;
        RECT 55.060 -58.080 56.240 -56.960 ;
        RECT 58.810 -58.080 59.990 -56.960 ;
        RECT 60.550 -57.220 61.720 -56.855 ;
        RECT 63.120 -57.220 64.290 -56.915 ;
        RECT 65.625 -57.220 66.795 -56.805 ;
        RECT 68.235 -57.220 69.405 -56.805 ;
        RECT 70.720 -57.220 71.890 -56.805 ;
        RECT 72.605 -57.220 73.375 -57.120 ;
        RECT 60.550 -57.520 73.375 -57.220 ;
        RECT 60.550 -57.985 61.720 -57.520 ;
        RECT 63.120 -58.045 64.290 -57.520 ;
        RECT 65.625 -57.935 66.795 -57.520 ;
        RECT 68.235 -57.935 69.405 -57.520 ;
        RECT 70.720 -57.935 71.890 -57.520 ;
        RECT 72.605 -57.850 73.375 -57.520 ;
        RECT 74.495 -58.120 75.665 -56.990 ;
        RECT 8.175 -65.165 9.345 -64.520 ;
        RECT 10.365 -65.165 10.665 -65.085 ;
        RECT 8.175 -65.465 10.665 -65.165 ;
        RECT 8.175 -65.650 9.345 -65.465 ;
        RECT 10.365 -66.730 10.665 -65.465 ;
        RECT 18.070 -65.650 19.240 -64.520 ;
        RECT 27.925 -65.650 29.095 -64.520 ;
        RECT 37.100 -65.650 38.270 -64.520 ;
        RECT 18.630 -66.730 18.930 -65.650 ;
        RECT 28.380 -66.730 28.680 -65.650 ;
        RECT 37.345 -66.730 37.645 -65.650 ;
        RECT 10.365 -67.030 37.645 -66.730 ;
        RECT 37.345 -75.015 37.645 -67.030 ;
        RECT 38.715 -72.170 39.015 -58.155 ;
        RECT 59.665 -68.805 60.835 -68.390 ;
        RECT 61.550 -68.805 62.720 -68.390 ;
        RECT 63.375 -68.805 64.545 -68.390 ;
        RECT 65.250 -68.805 66.420 -68.390 ;
        RECT 67.070 -68.805 68.240 -68.390 ;
        RECT 68.810 -68.805 69.980 -68.390 ;
        RECT 70.645 -68.805 71.815 -68.390 ;
        RECT 59.665 -69.105 71.815 -68.805 ;
        RECT 59.665 -69.520 60.835 -69.105 ;
        RECT 61.550 -69.520 62.720 -69.105 ;
        RECT 63.375 -69.520 64.545 -69.105 ;
        RECT 65.250 -69.520 66.420 -69.105 ;
        RECT 67.070 -69.520 68.240 -69.105 ;
        RECT 68.810 -69.520 69.980 -69.105 ;
        RECT 70.645 -69.520 71.815 -69.105 ;
        RECT 60.990 -70.195 62.160 -69.905 ;
        RECT 63.705 -70.195 64.005 -69.520 ;
        RECT 60.990 -70.495 64.900 -70.195 ;
        RECT 60.990 -71.035 62.160 -70.495 ;
        RECT 41.280 -72.170 42.050 -71.925 ;
        RECT 38.715 -72.470 42.050 -72.170 ;
        RECT 8.115 -75.430 9.285 -75.015 ;
        RECT 8.115 -75.730 11.090 -75.430 ;
        RECT 8.115 -76.145 9.285 -75.730 ;
        RECT 10.790 -77.095 11.090 -75.730 ;
        RECT 18.025 -76.145 19.195 -75.015 ;
        RECT 28.040 -76.145 29.210 -75.015 ;
        RECT 37.245 -76.145 38.415 -75.015 ;
        RECT 18.350 -77.095 18.650 -76.145 ;
        RECT 28.475 -77.095 28.775 -76.145 ;
        RECT 37.355 -77.095 37.655 -76.145 ;
        RECT 10.790 -77.395 37.955 -77.095 ;
        RECT 34.620 -77.845 34.920 -77.395 ;
        RECT 34.385 -78.575 35.155 -77.845 ;
        RECT 37.655 -84.000 37.955 -77.395 ;
        RECT 38.715 -80.125 39.015 -72.470 ;
        RECT 41.280 -72.655 42.050 -72.470 ;
        RECT 64.600 -78.405 64.900 -70.495 ;
        RECT 75.290 -70.830 75.590 -58.120 ;
        RECT 74.855 -71.960 76.025 -70.830 ;
        RECT 77.900 -71.960 79.070 -70.830 ;
        RECT 75.290 -74.475 75.590 -71.960 ;
        RECT 78.335 -72.425 78.635 -71.960 ;
        RECT 78.210 -73.145 78.990 -72.425 ;
        RECT 75.290 -74.775 77.995 -74.475 ;
        RECT 44.420 -79.535 45.590 -78.405 ;
        RECT 51.110 -79.535 52.280 -78.405 ;
        RECT 57.775 -79.535 58.945 -78.405 ;
        RECT 64.400 -79.535 65.570 -78.405 ;
        RECT 44.855 -80.125 45.155 -79.535 ;
        RECT 51.595 -80.125 51.895 -79.535 ;
        RECT 38.715 -80.425 51.895 -80.125 ;
        RECT 51.595 -82.365 51.895 -80.425 ;
        RECT 58.210 -80.135 58.510 -79.535 ;
        RECT 64.690 -80.135 64.990 -79.535 ;
        RECT 58.210 -80.435 64.990 -80.135 ;
        RECT 51.315 -83.095 52.085 -82.365 ;
        RECT 70.620 -82.800 71.790 -81.670 ;
        RECT 77.695 -81.685 77.995 -74.775 ;
        RECT 8.150 -85.130 9.320 -84.000 ;
        RECT 18.060 -85.130 19.230 -84.000 ;
        RECT 28.215 -85.130 29.385 -84.000 ;
        RECT 37.220 -85.130 38.390 -84.000 ;
        RECT 71.055 -84.675 71.355 -82.800 ;
        RECT 77.325 -82.815 78.495 -81.685 ;
        RECT 83.420 -82.780 84.590 -81.650 ;
        RECT 77.760 -83.790 78.060 -82.815 ;
        RECT 77.750 -84.675 78.060 -83.790 ;
        RECT 83.785 -83.745 84.085 -82.780 ;
        RECT 89.825 -82.825 90.995 -81.695 ;
        RECT 83.785 -84.045 84.105 -83.745 ;
        RECT 83.785 -84.675 84.085 -84.045 ;
        RECT 90.365 -84.675 90.665 -82.825 ;
        RECT 71.055 -84.975 90.665 -84.675 ;
        RECT 1.680 -86.800 1.995 -86.500 ;
        RECT 1.695 -87.850 1.995 -86.800 ;
        RECT 8.900 -87.850 9.200 -85.130 ;
        RECT 18.770 -87.850 19.070 -85.130 ;
        RECT 28.865 -85.795 29.165 -85.130 ;
        RECT 37.775 -85.795 38.075 -85.130 ;
        RECT 28.865 -86.095 38.075 -85.795 ;
        RECT 1.695 -88.150 19.070 -87.850 ;
        RECT 70.630 -91.610 71.800 -90.480 ;
        RECT 71.065 -92.360 71.365 -91.610 ;
        RECT 77.335 -91.960 78.505 -90.830 ;
        RECT 83.450 -91.960 84.620 -90.830 ;
        RECT 90.365 -91.820 90.665 -84.975 ;
        RECT 71.035 -93.700 71.365 -92.360 ;
        RECT 77.535 -93.700 77.835 -91.960 ;
        RECT 83.755 -93.700 84.055 -91.960 ;
        RECT 89.845 -92.950 91.015 -91.820 ;
        RECT 90.280 -93.700 90.580 -92.950 ;
        RECT 71.035 -94.000 90.580 -93.700 ;
      LAYER met4 ;
        RECT 49.475 -28.435 50.205 -27.705 ;
        RECT 75.770 -27.730 97.940 -6.625 ;
        RECT 75.590 -28.800 97.940 -27.730 ;
        RECT 55.085 -57.370 56.215 -56.955 ;
        RECT 58.835 -57.370 59.965 -56.955 ;
        RECT 55.085 -57.670 59.965 -57.370 ;
        RECT 55.085 -58.085 56.215 -57.670 ;
        RECT 58.120 -71.170 58.420 -57.670 ;
        RECT 58.835 -58.085 59.965 -57.670 ;
        RECT 58.120 -71.470 66.945 -71.170 ;
        RECT 66.645 -72.790 66.945 -71.470 ;
        RECT 66.645 -73.090 66.965 -72.790 ;
        RECT 66.665 -73.805 66.965 -73.090 ;
        RECT 78.235 -73.150 78.965 -72.420 ;
        RECT 78.450 -73.805 78.750 -73.150 ;
        RECT 66.665 -74.105 78.750 -73.805 ;
  END
END OpAmp
END LIBRARY

