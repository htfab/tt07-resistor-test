VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_WIDTH STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
  PROPERTY LEF58_SPACING "SPACING 1.27 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.84 ;" ;
END nwell

LAYER dnwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
  PROPERTY LEF58_ENCLOSURE "ENCLOSURE 0.4 LAYER nwell ;" ;
  PROPERTY LEF58_SPACING "SPACING 6.3 ;
  SPACING 4.5 LAYER nwell ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 3 ;" ;
END dnwell

LAYER diff
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.27 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.15 ;" ;
END diff

LAYER nsdm
  TYPE IMPLANT ;
  WIDTH 0.38 ;
  SPACING 0.38 ;
  AREA 0.265 ;
END nsdm

LAYER psdm
  TYPE IMPLANT ;
  WIDTH 0.38 ;
  SPACING 0.38 ;
  AREA 0.255 ;
END psdm

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER npc
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.27 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.27 ;" ;
END npc

LAYER licon
  TYPE CUT ;
  SPACING 0.17 ;
  WIDTH 0.17 ;
  ENCLOSURE BELOW 0.08 0.05 ;
  ENCLOSURE ABOVE 0.08 0.05 ;
  ANTENNAMODEL OXIDE1 ;
END licon

LAYER li
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.13 ;
  SPACING 0.17 ;
  RESISTANCE RPERSQ 12.2 ;
  CAPACITANCE CPERSQDIST 3.69e-05 ;
  THICKNESS 0.1 ;
  EDGECAPACITANCE 3.26e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 75 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 75 ) ( 0.0125 75 ) ( 0.0225 85.125 ) ( 22.5 10200 ) ) ;
END li

LAYER mcon
  TYPE CUT ;
  SPACING 0.19 ;
  WIDTH 0.17 ;
  ENCLOSURE ABOVE 0.06 0.03 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 3 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 3 ) ( 0.0125 3 ) ( 0.0225 3.405 ) ( 22.5 408 ) ) ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.14 ;
  OFFSET 0.185 0.185 ;
  AREA 0.083 ;
  SPACING 0.14 ;
  SPACING 0.28 RANGE 3.005 10000 ;
  SPACING 0.28 RANGE 3.005 10000 INFLUENCE 0.28 ;
  MINENCLOSEDAREA 0.14 ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 2.58e-05 ;
  THICKNESS 0.35 ;
  EDGECAPACITANCE 1.79e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met1

LAYER via1
  TYPE CUT ;
  SPACING 0.17 ;
  WIDTH 0.15 ;
  ENCLOSURE BELOW 0.085 0.055 ;
  ENCLOSURE ABOVE 0.085 0.055 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 6 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
END via1

LAYER met2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.14 ;
  OFFSET 0.185 0.185 ;
  AREA 0.0676 ;
  SPACING 0.14 ;
  SPACING 0.28 RANGE 3.005 10000 ;
  SPACING 0.28 RANGE 3.005 10000 INFLUENCE 0.28 ;
  MINENCLOSEDAREA 0.14 ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 1.75e-05 ;
  THICKNESS 0.35 ;
  EDGECAPACITANCE 1.22e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met2

LAYER via2
  TYPE CUT ;
  SPACING 0.2 ;
  WIDTH 0.2 ;
  ENCLOSURE BELOW 0.085 0.055 ;
  ENCLOSURE ABOVE 0.085 0.065 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 6 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.3 ;
  OFFSET 0.305 0.305 ;
  AREA 0.24 ;
  SPACING 0.3 ;
  SPACING 0.4 RANGE 3.005 10000 ;
  SPACING 0.4 RANGE 3.005 10000 INFLUENCE 0.4 ;
  RESISTANCE RPERSQ 0.047 ;
  CAPACITANCE CPERSQDIST 1.26e-05 ;
  THICKNESS 0.8 ;
  EDGECAPACITANCE 1.86e-06 ;
  ANTENNAMODEL OXIDE1 ;
END met3

LAYER via3
  TYPE CUT ;
  SPACING 0.2 ;
  WIDTH 0.2 ;
  ENCLOSURE BELOW 0.06 0.09 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 6 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.3 ;
  OFFSET 0.305 0.305 ;
  AREA 0.24 ;
  SPACING 0.3 ;
  SPACING 0.4 RANGE 3.005 10000 ;
  SPACING 0.4 RANGE 3.005 10000 INFLUENCE 0.4 ;
  RESISTANCE RPERSQ 0.047 ;
  CAPACITANCE CPERSQDIST 8.67e-06 ;
  THICKNESS 0.8 ;
  EDGECAPACITANCE 1.29e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met4

LAYER via4
  TYPE CUT ;
  SPACING 0.8 ;
  WIDTH 0.8 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 6 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.36 ;
  OFFSET 1.555 1.555 ;
  SPACING 0.36 ;
  RESISTANCE RPERSQ 0.0285 ;
  CAPACITANCE CPERSQDIST 6.48e-06 ;
  THICKNESS 1.2 ;
  EDGECAPACITANCE 4.96e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met5

LAYER rdl
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 10 ;
  SPACING 10 ;
  RESISTANCE RPERSQ 0.005 ;
  CAPACITANCE CPERSQDIST 2.66e-06 ;
  THICKNESS 2 ;
  EDGECAPACITANCE 6.2e-06 ;
  ANTENNAMODEL OXIDE1 ;
END rdl

VIARULE M4M5 GENERATE DEFAULT
  LAYER met5 ;
    ENCLOSURE 0.31 0.31 ;
  LAYER met4 ;
    ENCLOSURE 0.19 0.19 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.6 BY 1.6 ;
    RESISTANCE 0.380000 ;
END M4M5

VIARULE M3M4 GENERATE DEFAULT
  LAYER met4 ;
    ENCLOSURE 0.065 0.065 ;
  LAYER met3 ;
    ENCLOSURE 0.09 0.06 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
    RESISTANCE 3.410000 ;
END M3M4

VIARULE M2M3 GENERATE DEFAULT
  LAYER met3 ;
    ENCLOSURE 0.065 0.065 ;
  LAYER met2 ;
    ENCLOSURE 0.085 0.065 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
    RESISTANCE 3.410000 ;
END M2M3

VIARULE M1M2 GENERATE DEFAULT
  LAYER met2 ;
    ENCLOSURE 0.085 0.055 ;
  LAYER met1 ;
    ENCLOSURE 0.085 0.055 ;
  LAYER via1 ;
    RECT -0.075 -0.075 0.075 0.075 ;
    SPACING 0.32 BY 0.32 ;
    RESISTANCE 4.500000 ;
END M1M2

VIARULE L1M1 GENERATE
  LAYER met1 ;
    ENCLOSURE 0.06 0.03 ;
  LAYER li ;
    ENCLOSURE 0 0 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
    SPACING 0.36 BY 0.36 ;
    RESISTANCE 9.300000 ;
END L1M1

VIARULE PYL1 GENERATE
  LAYER poly ;
    ENCLOSURE 0.08 0.05 ;
  LAYER li ;
    ENCLOSURE 0.08 0 ;
  LAYER licon ;
    RECT -0.085 -0.085 0.085 0.085 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 145.279999 ;
END PYL1

VIARULE DFL1 GENERATE
  LAYER li ;
    ENCLOSURE 0.08 0.08 ;
  LAYER diff ;
    ENCLOSURE 0.12 0.12 ;
  LAYER licon ;
    RECT -0.085 -0.085 0.085 0.085 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 600.000000 ;
END DFL1

VIARULE NPDF GENERATE
  LAYER li ;
    ENCLOSURE 0.08 0.08 ;
  LAYER diff ;
    ENCLOSURE 0.12 0.12 ;
  LAYER licon ;
    RECT -0.085 -0.085 0.085 0.085 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 600.000000 ;
END NPDF

VIARULE PPDF GENERATE
  LAYER li ;
    ENCLOSURE 0.08 0.08 ;
  LAYER diff ;
    ENCLOSURE 0.12 0.12 ;
  LAYER licon ;
    RECT -0.085 -0.085 0.085 0.085 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 600.000000 ;
END PPDF

VIARULE NTAP GENERATE
  LAYER li ;
    ENCLOSURE 0.08 0.08 ;
  LAYER diff ;
    ENCLOSURE 0.12 0.12 ;
  LAYER licon ;
    RECT -0.085 -0.085 0.085 0.085 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 600.000000 ;
END NTAP

VIARULE PTAP GENERATE
  LAYER li ;
    ENCLOSURE 0.08 0.08 ;
  LAYER diff ;
    ENCLOSURE 0.12 0.12 ;
  LAYER licon ;
    RECT -0.085 -0.085 0.085 0.085 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 600.000000 ;
END PTAP

MACRO tt_um_resistor_davidparent
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.8 221.84 36.315 223.575 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.08 222.28 2.385 223.435 ;
    END
  END VPWR
END tt_um_resistor_davidparent

END LIBRARY
