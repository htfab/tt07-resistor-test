VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Burrows_Katie
  CLASS BLOCK ;
  FOREIGN tt_um_Burrows_Katie ;
  ORIGIN -54.365 -35.020 ;
  SIZE 158.355 BY 225.760 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 57.065 54.275 57.075 54.285 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 211.645 43.985 211.655 43.995 ;
    END
  END VPWR
  OBS
      LAYER pwell ;
        RECT 105.010 247.200 105.680 247.280 ;
        RECT 105.010 244.410 110.950 247.200 ;
      LAYER nwell ;
        RECT 150.485 245.390 156.905 250.670 ;
        RECT 158.565 245.390 164.985 250.670 ;
      LAYER pwell ;
        RECT 105.010 244.330 105.680 244.410 ;
        RECT 105.010 242.500 105.680 242.580 ;
        RECT 105.010 239.710 110.950 242.500 ;
      LAYER nwell ;
        RECT 115.670 241.320 118.090 244.600 ;
        RECT 144.650 241.355 147.070 244.635 ;
      LAYER pwell ;
        RECT 105.010 239.630 105.680 239.710 ;
      LAYER nwell ;
        RECT 150.485 238.400 156.905 243.680 ;
        RECT 158.565 238.400 164.985 243.680 ;
      LAYER pwell ;
        RECT 105.010 235.965 105.680 236.045 ;
        RECT 105.010 233.175 110.950 235.965 ;
        RECT 105.010 233.095 105.680 233.175 ;
      LAYER nwell ;
        RECT 129.195 232.010 135.615 237.290 ;
        RECT 150.485 231.410 156.905 236.690 ;
        RECT 158.565 231.410 164.985 236.690 ;
      LAYER pwell ;
        RECT 105.010 231.155 105.680 231.235 ;
        RECT 105.010 228.365 110.950 231.155 ;
        RECT 105.010 228.285 105.680 228.365 ;
      LAYER nwell ;
        RECT 129.195 225.095 135.615 230.375 ;
        RECT 150.485 224.385 156.905 229.665 ;
        RECT 158.565 224.385 164.985 229.665 ;
      LAYER pwell ;
        RECT 97.915 222.760 98.585 222.840 ;
        RECT 97.915 219.970 105.855 222.760 ;
        RECT 97.915 219.890 98.585 219.970 ;
        RECT 97.915 218.285 98.585 218.365 ;
        RECT 97.915 215.495 105.855 218.285 ;
        RECT 97.915 215.415 98.585 215.495 ;
        RECT 97.915 213.670 98.585 213.750 ;
        RECT 97.915 210.880 105.855 213.670 ;
        RECT 97.915 210.800 98.585 210.880 ;
        RECT 97.895 208.095 98.565 208.175 ;
        RECT 97.895 205.305 105.835 208.095 ;
      LAYER nwell ;
        RECT 141.045 207.385 143.465 210.665 ;
        RECT 158.790 205.770 165.210 211.050 ;
      LAYER pwell ;
        RECT 97.895 205.225 98.565 205.305 ;
        RECT 97.895 203.580 98.565 203.660 ;
        RECT 97.895 200.790 105.835 203.580 ;
        RECT 97.895 200.710 98.565 200.790 ;
        RECT 97.895 198.990 98.565 199.070 ;
        RECT 97.895 196.200 105.835 198.990 ;
      LAYER nwell ;
        RECT 141.040 197.385 143.460 200.665 ;
        RECT 158.790 198.660 165.210 203.940 ;
      LAYER pwell ;
        RECT 97.895 196.120 98.565 196.200 ;
        RECT 95.795 142.245 96.465 142.325 ;
        RECT 95.795 137.455 101.735 142.245 ;
        RECT 95.795 137.375 96.465 137.455 ;
      LAYER nwell ;
        RECT 105.060 137.265 111.480 142.545 ;
        RECT 115.210 137.265 121.630 142.545 ;
        RECT 124.490 137.220 130.910 142.500 ;
      LAYER pwell ;
        RECT 95.795 132.430 96.465 132.510 ;
        RECT 95.795 127.640 101.735 132.430 ;
        RECT 95.795 127.560 96.465 127.640 ;
      LAYER nwell ;
        RECT 105.060 127.370 111.480 132.650 ;
        RECT 115.210 127.390 121.630 132.670 ;
        RECT 124.490 127.330 130.910 132.610 ;
      LAYER pwell ;
        RECT 95.795 122.270 96.465 122.350 ;
        RECT 95.795 117.480 101.735 122.270 ;
        RECT 95.795 117.400 96.465 117.480 ;
      LAYER nwell ;
        RECT 105.060 117.325 111.480 122.605 ;
        RECT 115.210 117.450 121.630 122.730 ;
        RECT 124.445 117.495 130.865 122.775 ;
        RECT 147.890 116.235 154.310 129.205 ;
        RECT 166.235 116.235 172.655 129.205 ;
      LAYER pwell ;
        RECT 95.795 113.205 96.465 113.285 ;
        RECT 95.795 108.415 101.735 113.205 ;
        RECT 95.795 108.335 96.465 108.415 ;
      LAYER nwell ;
        RECT 105.060 108.125 111.480 113.405 ;
        RECT 115.210 108.030 121.630 113.310 ;
        RECT 124.490 107.935 130.910 113.215 ;
      LAYER pwell ;
        RECT 101.480 104.990 102.150 105.070 ;
        RECT 101.480 101.200 108.420 104.990 ;
        RECT 101.480 101.120 102.150 101.200 ;
        RECT 101.480 98.300 102.150 98.380 ;
        RECT 101.480 94.510 108.420 98.300 ;
        RECT 101.480 94.430 102.150 94.510 ;
        RECT 101.480 91.610 102.150 91.690 ;
        RECT 101.480 87.820 108.420 91.610 ;
      LAYER nwell ;
        RECT 114.405 89.470 122.825 103.210 ;
        RECT 126.760 89.890 135.180 103.690 ;
        RECT 147.585 97.945 154.005 110.915 ;
        RECT 166.240 97.700 172.660 110.670 ;
      LAYER pwell ;
        RECT 101.480 87.740 102.150 87.820 ;
        RECT 101.480 84.970 102.150 85.050 ;
        RECT 101.480 81.180 108.420 84.970 ;
        RECT 101.480 81.100 102.150 81.180 ;
        RECT 88.010 78.770 88.680 78.850 ;
        RECT 98.135 78.770 98.805 78.850 ;
        RECT 88.010 74.980 95.050 78.770 ;
        RECT 98.135 74.980 105.175 78.770 ;
        RECT 88.010 74.900 88.680 74.980 ;
        RECT 98.135 74.900 98.805 74.980 ;
      LAYER nwell ;
        RECT 114.660 72.765 123.080 86.505 ;
        RECT 126.780 72.245 135.200 86.045 ;
        RECT 163.425 78.670 171.845 91.010 ;
      LAYER pwell ;
        RECT 88.010 72.075 88.680 72.155 ;
        RECT 98.135 72.075 98.805 72.155 ;
        RECT 88.010 68.285 95.050 72.075 ;
        RECT 98.135 68.285 105.175 72.075 ;
        RECT 122.490 69.315 123.160 69.395 ;
        RECT 109.040 69.140 109.710 69.220 ;
        RECT 88.010 68.205 88.680 68.285 ;
        RECT 98.135 68.205 98.805 68.285 ;
        RECT 109.040 67.720 116.980 69.140 ;
        RECT 122.490 67.895 130.430 69.315 ;
        RECT 122.490 67.815 123.160 67.895 ;
        RECT 109.040 67.640 109.710 67.720 ;
        RECT 88.010 65.960 88.680 66.040 ;
        RECT 98.135 65.960 98.805 66.040 ;
        RECT 88.010 62.170 95.050 65.960 ;
        RECT 98.135 62.170 105.175 65.960 ;
        RECT 88.010 62.090 88.680 62.170 ;
        RECT 98.135 62.090 98.805 62.170 ;
        RECT 88.010 59.555 88.680 59.635 ;
        RECT 98.135 59.555 98.805 59.635 ;
        RECT 88.010 55.765 95.050 59.555 ;
        RECT 98.135 55.765 105.175 59.555 ;
        RECT 88.010 55.685 88.680 55.765 ;
        RECT 98.135 55.685 98.805 55.765 ;
      LAYER li1 ;
        RECT 151.360 250.650 151.890 251.180 ;
        RECT 159.640 250.650 160.170 251.180 ;
        RECT 151.475 250.255 151.775 250.650 ;
        RECT 151.170 250.085 155.920 250.255 ;
        RECT 156.355 249.590 156.685 250.335 ;
        RECT 159.755 250.255 160.055 250.650 ;
        RECT 159.250 250.085 164.000 250.255 ;
        RECT 156.970 249.590 157.500 249.725 ;
        RECT 156.355 249.260 157.500 249.590 ;
        RECT 105.180 246.285 105.510 247.110 ;
        RECT 106.215 247.030 106.915 248.220 ;
        RECT 149.965 247.990 150.565 248.590 ;
        RECT 105.945 246.860 110.695 247.030 ;
        RECT 104.270 245.585 105.510 246.285 ;
        RECT 105.180 244.500 105.510 245.585 ;
        RECT 111.375 245.440 111.905 245.970 ;
        RECT 151.170 245.805 155.920 245.975 ;
        RECT 155.605 245.390 155.775 245.805 ;
        RECT 156.355 245.725 156.685 249.260 ;
        RECT 156.970 249.195 157.500 249.260 ;
        RECT 164.435 249.435 164.765 250.335 ;
        RECT 165.070 249.435 165.600 249.575 ;
        RECT 164.435 249.105 165.600 249.435 ;
        RECT 158.160 248.130 158.760 248.730 ;
        RECT 159.250 245.805 164.000 245.975 ;
        RECT 159.455 245.660 159.760 245.805 ;
        RECT 164.435 245.725 164.765 249.105 ;
        RECT 165.070 249.045 165.600 249.105 ;
        RECT 159.460 245.390 159.760 245.660 ;
        RECT 105.945 244.580 110.695 244.750 ;
        RECT 116.475 244.650 117.005 245.180 ;
        RECT 145.560 244.650 146.090 245.180 ;
        RECT 155.425 244.860 155.955 245.390 ;
        RECT 159.345 244.860 159.875 245.390 ;
        RECT 106.015 244.250 106.315 244.580 ;
        RECT 105.900 243.720 106.430 244.250 ;
        RECT 116.590 244.185 116.760 244.650 ;
        RECT 117.560 244.265 117.890 244.285 ;
        RECT 116.395 244.015 117.065 244.185 ;
        RECT 105.180 241.385 105.510 242.410 ;
        RECT 106.205 242.330 106.905 243.155 ;
        RECT 114.935 242.940 115.825 243.830 ;
        RECT 105.945 242.160 110.695 242.330 ;
        RECT 116.395 241.840 117.065 241.905 ;
        RECT 104.270 240.685 105.510 241.385 ;
        RECT 116.380 241.735 117.065 241.840 ;
        RECT 116.380 241.375 116.780 241.735 ;
        RECT 117.540 241.655 117.890 244.265 ;
        RECT 145.685 244.220 145.985 244.650 ;
        RECT 145.375 244.050 146.045 244.220 ;
        RECT 145.685 244.015 145.985 244.050 ;
        RECT 143.845 242.940 144.735 243.830 ;
        RECT 145.375 241.770 146.045 241.940 ;
        RECT 146.520 241.830 146.850 244.300 ;
        RECT 151.360 243.455 151.890 243.985 ;
        RECT 159.640 243.455 160.170 243.985 ;
        RECT 151.475 243.265 151.775 243.455 ;
        RECT 151.170 243.095 155.920 243.265 ;
        RECT 111.375 240.785 111.905 241.315 ;
        RECT 116.295 240.845 116.825 241.375 ;
        RECT 105.180 239.800 105.510 240.685 ;
        RECT 117.560 240.300 117.890 241.655 ;
        RECT 145.685 241.395 145.985 241.770 ;
        RECT 146.495 241.690 146.850 241.830 ;
        RECT 156.355 242.670 156.685 243.345 ;
        RECT 159.755 243.265 160.055 243.455 ;
        RECT 159.250 243.095 164.000 243.265 ;
        RECT 156.990 242.670 157.520 242.810 ;
        RECT 156.355 242.340 157.520 242.670 ;
        RECT 145.560 240.865 146.090 241.395 ;
        RECT 146.495 240.395 146.825 241.690 ;
        RECT 149.965 240.815 150.565 241.415 ;
        RECT 105.945 239.880 110.695 240.050 ;
        RECT 105.975 239.440 106.275 239.880 ;
        RECT 117.560 239.870 118.100 240.300 ;
        RECT 117.570 239.770 118.100 239.870 ;
        RECT 146.370 239.865 146.900 240.395 ;
        RECT 105.860 238.910 106.390 239.440 ;
        RECT 151.170 238.815 155.920 238.985 ;
        RECT 155.690 238.325 155.860 238.815 ;
        RECT 156.355 238.735 156.685 242.340 ;
        RECT 156.990 242.280 157.520 242.340 ;
        RECT 164.435 242.670 164.765 243.345 ;
        RECT 165.070 242.670 165.600 242.810 ;
        RECT 164.435 242.340 165.600 242.670 ;
        RECT 158.160 241.050 158.760 241.650 ;
        RECT 159.250 238.815 164.000 238.985 ;
        RECT 159.545 238.325 159.845 238.815 ;
        RECT 164.435 238.735 164.765 242.340 ;
        RECT 165.070 242.280 165.600 242.340 ;
        RECT 133.840 236.875 134.540 238.095 ;
        RECT 155.510 237.795 156.040 238.325 ;
        RECT 159.430 237.795 159.960 238.325 ;
        RECT 105.180 234.850 105.510 235.875 ;
        RECT 106.130 235.795 106.830 236.725 ;
        RECT 129.880 236.705 134.630 236.875 ;
        RECT 135.065 236.835 135.395 236.955 ;
        RECT 135.065 236.135 136.365 236.835 ;
        RECT 151.360 236.480 151.890 237.010 ;
        RECT 159.640 236.550 160.170 237.080 ;
        RECT 151.475 236.275 151.775 236.480 ;
        RECT 105.945 235.625 110.695 235.795 ;
        RECT 104.270 234.150 105.510 234.850 ;
        RECT 111.375 234.390 111.905 234.920 ;
        RECT 128.640 234.405 129.170 234.935 ;
        RECT 105.180 233.265 105.510 234.150 ;
        RECT 105.945 233.345 110.695 233.515 ;
        RECT 106.030 233.020 106.330 233.345 ;
        RECT 105.915 232.490 106.445 233.020 ;
        RECT 129.880 232.425 134.630 232.595 ;
        RECT 130.200 232.040 130.500 232.425 ;
        RECT 135.065 232.345 135.395 236.135 ;
        RECT 151.170 236.105 155.920 236.275 ;
        RECT 156.355 235.495 156.685 236.355 ;
        RECT 159.755 236.275 160.055 236.550 ;
        RECT 159.250 236.105 164.000 236.275 ;
        RECT 156.990 235.495 157.520 235.700 ;
        RECT 156.355 235.170 157.520 235.495 ;
        RECT 164.435 235.495 164.765 236.355 ;
        RECT 165.070 235.495 165.600 235.700 ;
        RECT 164.435 235.170 165.600 235.495 ;
        RECT 156.355 235.165 157.420 235.170 ;
        RECT 164.435 235.165 165.500 235.170 ;
        RECT 149.965 233.865 150.565 234.465 ;
        RECT 105.180 230.160 105.510 231.065 ;
        RECT 106.185 230.985 106.885 231.800 ;
        RECT 130.085 231.510 130.615 232.040 ;
        RECT 151.170 231.825 155.920 231.995 ;
        RECT 155.690 231.445 155.860 231.825 ;
        RECT 156.355 231.745 156.685 235.165 ;
        RECT 158.160 234.180 158.760 234.780 ;
        RECT 159.250 231.825 164.000 231.995 ;
        RECT 159.545 231.445 159.845 231.825 ;
        RECT 164.435 231.745 164.765 235.165 ;
        RECT 105.945 230.815 110.695 230.985 ;
        RECT 104.270 229.460 105.510 230.160 ;
        RECT 133.840 229.960 134.540 230.990 ;
        RECT 155.510 230.915 156.040 231.445 ;
        RECT 159.430 230.915 159.960 231.445 ;
        RECT 105.180 228.455 105.510 229.460 ;
        RECT 111.375 229.345 111.905 229.875 ;
        RECT 129.880 229.790 134.630 229.960 ;
        RECT 135.065 229.940 135.395 230.040 ;
        RECT 135.065 229.240 136.365 229.940 ;
        RECT 151.360 229.505 151.890 230.035 ;
        RECT 159.640 229.570 160.170 230.100 ;
        RECT 151.540 229.250 151.710 229.505 ;
        RECT 105.945 228.535 110.695 228.705 ;
        RECT 105.995 228.200 106.295 228.535 ;
        RECT 105.915 227.670 106.445 228.200 ;
        RECT 128.620 227.130 129.150 227.660 ;
        RECT 129.880 225.510 134.630 225.680 ;
        RECT 130.200 225.175 130.500 225.510 ;
        RECT 135.065 225.430 135.395 229.240 ;
        RECT 151.170 229.080 155.920 229.250 ;
        RECT 156.355 228.395 156.685 229.330 ;
        RECT 159.755 229.250 160.055 229.570 ;
        RECT 159.250 229.080 164.000 229.250 ;
        RECT 156.990 228.395 157.520 228.635 ;
        RECT 156.355 228.105 157.520 228.395 ;
        RECT 156.355 228.065 157.420 228.105 ;
        RECT 149.965 226.840 150.565 227.440 ;
        RECT 130.085 224.645 130.615 225.175 ;
        RECT 151.170 224.800 155.920 224.970 ;
        RECT 155.690 224.285 155.860 224.800 ;
        RECT 156.355 224.720 156.685 228.065 ;
        RECT 164.435 227.955 164.765 229.330 ;
        RECT 165.070 227.955 165.600 228.195 ;
        RECT 164.435 227.665 165.600 227.955 ;
        RECT 164.435 227.625 165.500 227.665 ;
        RECT 158.160 226.840 158.760 227.440 ;
        RECT 159.250 224.800 164.000 224.970 ;
        RECT 159.545 224.285 159.845 224.800 ;
        RECT 164.435 224.720 164.765 227.625 ;
        RECT 98.085 222.590 98.415 222.670 ;
        RECT 98.950 222.590 99.650 223.765 ;
        RECT 155.510 223.755 156.040 224.285 ;
        RECT 159.430 223.755 159.960 224.285 ;
        RECT 97.025 221.890 98.415 222.590 ;
        RECT 98.830 222.420 105.620 222.590 ;
        RECT 98.085 220.060 98.415 221.890 ;
        RECT 106.235 221.075 106.765 221.605 ;
        RECT 98.830 220.140 105.620 220.310 ;
        RECT 105.315 219.780 105.615 220.140 ;
        RECT 105.225 219.250 105.755 219.780 ;
        RECT 110.920 219.060 111.090 220.940 ;
        RECT 171.255 220.270 171.425 220.940 ;
        RECT 98.085 218.135 98.415 218.195 ;
        RECT 97.025 217.435 98.415 218.135 ;
        RECT 98.950 218.115 99.650 219.035 ;
        RECT 98.830 217.945 105.620 218.115 ;
        RECT 98.085 215.585 98.415 217.435 ;
        RECT 106.235 216.620 106.765 217.150 ;
        RECT 110.920 216.640 111.090 218.520 ;
        RECT 171.255 217.850 171.425 219.730 ;
        RECT 98.830 215.665 105.620 215.835 ;
        RECT 105.310 215.265 105.610 215.665 ;
        RECT 105.225 214.735 105.755 215.265 ;
        RECT 98.085 213.535 98.415 213.580 ;
        RECT 97.025 212.835 98.415 213.535 ;
        RECT 98.950 213.500 99.650 214.470 ;
        RECT 110.920 214.220 111.090 216.100 ;
        RECT 171.255 215.430 171.425 217.310 ;
        RECT 171.255 214.220 171.425 214.890 ;
        RECT 98.830 213.330 105.620 213.500 ;
        RECT 98.085 210.970 98.415 212.835 ;
        RECT 106.235 211.925 106.765 212.455 ;
        RECT 98.830 211.050 105.620 211.220 ;
        RECT 105.315 210.665 105.615 211.050 ;
        RECT 105.225 210.135 105.755 210.665 ;
        RECT 141.625 210.635 142.155 211.165 ;
        RECT 159.375 210.635 160.075 211.655 ;
        RECT 141.770 210.250 142.070 210.635 ;
        RECT 159.375 210.530 164.225 210.635 ;
        RECT 159.475 210.465 164.225 210.530 ;
        RECT 141.770 210.080 142.440 210.250 ;
        RECT 141.770 210.020 142.070 210.080 ;
        RECT 98.065 207.990 98.395 208.005 ;
        RECT 97.025 207.290 98.395 207.990 ;
        RECT 98.865 207.925 99.565 208.900 ;
        RECT 140.270 208.630 141.160 209.520 ;
        RECT 142.915 209.275 143.245 210.330 ;
        RECT 164.660 209.975 164.990 210.715 ;
        RECT 164.660 209.275 166.105 209.975 ;
        RECT 142.915 208.575 144.180 209.275 ;
        RECT 98.810 207.755 105.600 207.925 ;
        RECT 141.770 207.800 142.440 207.970 ;
        RECT 98.065 205.395 98.395 207.290 ;
        RECT 141.770 207.195 142.070 207.800 ;
        RECT 142.915 207.720 143.245 208.575 ;
        RECT 158.130 207.775 158.730 208.375 ;
        RECT 106.210 206.215 106.740 206.745 ;
        RECT 141.650 206.665 142.180 207.195 ;
        RECT 159.575 206.355 160.275 206.365 ;
        RECT 159.475 206.185 164.225 206.355 ;
        RECT 98.810 205.475 105.600 205.645 ;
        RECT 98.065 203.350 98.395 203.490 ;
        RECT 98.865 203.410 99.565 204.450 ;
        RECT 104.880 204.440 105.580 205.475 ;
        RECT 159.575 205.240 160.275 206.185 ;
        RECT 164.660 206.105 164.990 209.275 ;
        RECT 159.375 203.525 160.075 204.485 ;
        RECT 159.375 203.435 164.225 203.525 ;
        RECT 97.090 202.650 98.395 203.350 ;
        RECT 98.810 203.240 105.600 203.410 ;
        RECT 159.475 203.355 164.225 203.435 ;
        RECT 164.660 203.420 164.990 203.605 ;
        RECT 98.065 200.880 98.395 202.650 ;
        RECT 164.660 202.720 166.015 203.420 ;
        RECT 106.240 201.905 106.770 202.435 ;
        RECT 98.810 200.960 105.600 201.130 ;
        RECT 104.880 199.900 105.580 200.960 ;
        RECT 141.640 200.575 142.170 201.105 ;
        RECT 146.365 200.605 146.895 201.135 ;
        RECT 158.130 200.985 158.730 201.585 ;
        RECT 141.775 200.250 142.075 200.575 ;
        RECT 141.765 200.080 142.435 200.250 ;
        RECT 141.775 200.010 142.075 200.080 ;
        RECT 98.065 198.885 98.395 198.900 ;
        RECT 97.025 198.185 98.395 198.885 ;
        RECT 98.865 198.820 99.565 199.875 ;
        RECT 98.810 198.650 105.600 198.820 ;
        RECT 140.360 198.670 141.250 199.560 ;
        RECT 142.910 199.320 143.240 200.330 ;
        RECT 98.065 196.290 98.395 198.185 ;
        RECT 142.910 198.620 144.245 199.320 ;
        RECT 159.475 199.075 164.225 199.245 ;
        RECT 106.220 197.305 106.750 197.835 ;
        RECT 141.765 197.800 142.435 197.970 ;
        RECT 141.775 197.205 142.075 197.800 ;
        RECT 142.910 197.720 143.240 198.620 ;
        RECT 159.575 198.100 160.275 199.075 ;
        RECT 164.660 198.995 164.990 202.720 ;
        RECT 141.650 196.675 142.180 197.205 ;
        RECT 98.810 196.370 105.600 196.540 ;
        RECT 104.860 195.150 105.560 196.370 ;
        RECT 98.280 191.400 98.450 193.280 ;
        RECT 163.285 192.610 163.455 193.280 ;
        RECT 98.280 188.980 98.450 190.860 ;
        RECT 163.285 190.190 163.455 192.070 ;
        RECT 98.280 186.560 98.450 188.440 ;
        RECT 163.285 187.770 163.455 189.650 ;
        RECT 98.280 184.140 98.450 186.020 ;
        RECT 163.285 185.350 163.455 187.230 ;
        RECT 98.280 181.720 98.450 183.600 ;
        RECT 163.285 182.930 163.455 184.810 ;
        RECT 98.280 179.300 98.450 181.180 ;
        RECT 163.285 180.510 163.455 182.390 ;
        RECT 98.280 176.880 98.450 178.760 ;
        RECT 163.285 178.090 163.455 179.970 ;
        RECT 98.280 174.460 98.450 176.340 ;
        RECT 163.285 175.670 163.455 177.550 ;
        RECT 163.285 174.460 163.455 175.130 ;
        RECT 96.600 142.755 97.130 142.925 ;
        RECT 105.585 142.765 106.115 142.935 ;
        RECT 115.820 142.765 116.350 142.935 ;
        RECT 95.965 140.910 96.295 142.155 ;
        RECT 96.775 142.075 96.945 142.755 ;
        RECT 105.760 142.130 105.930 142.765 ;
        RECT 96.730 141.905 101.480 142.075 ;
        RECT 105.745 141.960 110.495 142.130 ;
        RECT 96.775 141.900 96.945 141.905 ;
        RECT 94.610 139.910 96.295 140.910 ;
        RECT 110.930 140.335 111.260 142.210 ;
        RECT 115.995 142.130 116.165 142.765 ;
        RECT 115.895 141.960 120.645 142.130 ;
        RECT 121.080 140.375 121.410 142.210 ;
        RECT 129.210 142.085 129.910 143.515 ;
        RECT 125.175 141.915 129.925 142.085 ;
        RECT 129.210 141.905 129.910 141.915 ;
        RECT 95.965 137.545 96.295 139.910 ;
        RECT 102.140 139.770 102.670 140.300 ;
        RECT 110.930 140.265 112.305 140.335 ;
        RECT 121.080 140.265 122.515 140.375 ;
        RECT 110.930 140.095 112.590 140.265 ;
        RECT 121.080 140.095 122.615 140.265 ;
        RECT 110.930 140.005 112.305 140.095 ;
        RECT 121.080 140.045 122.515 140.095 ;
        RECT 104.580 137.805 105.110 138.335 ;
        RECT 96.730 137.625 101.480 137.795 ;
        RECT 105.745 137.680 110.495 137.850 ;
        RECT 96.800 137.175 96.970 137.625 ;
        RECT 105.785 137.210 105.955 137.680 ;
        RECT 110.930 137.600 111.260 140.005 ;
        RECT 114.740 137.775 115.270 138.305 ;
        RECT 115.895 137.680 120.645 137.850 ;
        RECT 96.340 136.175 97.340 137.175 ;
        RECT 105.325 136.210 106.325 137.210 ;
        RECT 116.280 137.150 116.450 137.680 ;
        RECT 121.080 137.600 121.410 140.045 ;
        RECT 123.940 139.565 124.470 140.095 ;
        RECT 125.175 137.635 129.925 137.805 ;
        RECT 115.820 136.150 116.820 137.150 ;
        RECT 125.195 137.130 125.365 137.635 ;
        RECT 124.790 136.240 125.680 137.130 ;
        RECT 130.360 136.595 130.690 142.165 ;
        RECT 133.515 138.270 133.685 138.940 ;
        RECT 130.075 136.550 130.690 136.595 ;
        RECT 129.975 136.380 130.690 136.550 ;
        RECT 130.075 136.265 130.690 136.380 ;
        RECT 133.515 135.850 133.685 137.730 ;
        RECT 174.350 137.060 174.520 138.940 ;
        RECT 96.600 133.905 97.130 134.075 ;
        RECT 95.965 131.115 96.295 132.340 ;
        RECT 96.775 132.260 96.945 133.905 ;
        RECT 105.585 132.805 106.115 132.975 ;
        RECT 115.820 132.825 116.350 132.995 ;
        RECT 96.730 132.090 101.480 132.260 ;
        RECT 105.760 132.235 105.930 132.805 ;
        RECT 105.745 132.065 110.495 132.235 ;
        RECT 94.610 130.115 96.295 131.115 ;
        RECT 95.965 127.730 96.295 130.115 ;
        RECT 102.160 129.660 102.690 130.190 ;
        RECT 110.930 129.945 111.260 132.315 ;
        RECT 115.995 132.255 116.165 132.825 ;
        RECT 114.740 131.580 115.270 132.110 ;
        RECT 115.895 132.085 120.645 132.255 ;
        RECT 121.080 130.050 121.410 132.335 ;
        RECT 129.210 132.195 129.910 133.610 ;
        RECT 133.515 133.430 133.685 135.310 ;
        RECT 174.350 134.640 174.520 136.520 ;
        RECT 174.350 133.430 174.520 134.100 ;
        RECT 125.175 132.025 129.925 132.195 ;
        RECT 129.210 132.000 129.910 132.025 ;
        RECT 110.930 129.915 112.350 129.945 ;
        RECT 121.080 129.915 122.515 130.050 ;
        RECT 110.930 129.745 112.590 129.915 ;
        RECT 121.080 129.745 122.615 129.915 ;
        RECT 110.930 129.615 112.350 129.745 ;
        RECT 121.080 129.720 122.515 129.745 ;
        RECT 96.730 127.810 101.480 127.980 ;
        RECT 104.580 127.875 105.110 128.405 ;
        RECT 96.800 127.265 96.970 127.810 ;
        RECT 105.745 127.785 110.495 127.955 ;
        RECT 105.785 127.300 105.955 127.785 ;
        RECT 110.930 127.705 111.260 129.615 ;
        RECT 115.895 127.805 120.645 127.975 ;
        RECT 96.340 126.265 97.340 127.265 ;
        RECT 105.325 126.300 106.325 127.300 ;
        RECT 116.280 127.255 116.450 127.805 ;
        RECT 121.080 127.725 121.410 129.720 ;
        RECT 123.960 129.600 124.490 130.130 ;
        RECT 125.175 127.745 129.925 127.915 ;
        RECT 115.820 126.255 116.820 127.255 ;
        RECT 125.195 127.230 125.365 127.745 ;
        RECT 124.790 126.340 125.680 127.230 ;
        RECT 130.360 127.080 130.690 132.275 ;
        RECT 143.805 129.540 144.335 130.070 ;
        RECT 147.010 129.475 148.010 130.475 ;
        RECT 162.840 130.135 163.370 130.665 ;
        RECT 148.700 129.695 149.230 129.865 ;
        RECT 145.105 127.775 146.105 128.750 ;
        RECT 146.770 128.590 147.300 128.615 ;
        RECT 146.770 128.445 147.385 128.590 ;
        RECT 147.140 128.420 147.385 128.445 ;
        RECT 145.105 127.750 146.945 127.775 ;
        RECT 145.680 127.605 146.945 127.750 ;
        RECT 130.075 127.030 130.690 127.080 ;
        RECT 129.975 126.860 130.690 127.030 ;
        RECT 130.075 126.750 130.690 126.860 ;
        RECT 144.075 126.185 145.075 127.185 ;
        RECT 146.775 127.115 146.945 127.605 ;
        RECT 147.215 127.530 147.385 128.420 ;
        RECT 147.735 128.150 147.905 129.475 ;
        RECT 148.880 128.790 149.050 129.695 ;
        RECT 165.340 129.475 166.340 130.475 ;
        RECT 167.030 129.695 167.560 129.865 ;
        RECT 148.575 128.620 153.325 128.790 ;
        RECT 148.575 128.150 153.325 128.160 ;
        RECT 147.735 127.990 153.325 128.150 ;
        RECT 147.735 127.980 148.705 127.990 ;
        RECT 153.760 127.625 154.090 128.870 ;
        RECT 155.140 127.625 156.140 128.065 ;
        RECT 163.435 127.775 164.435 128.750 ;
        RECT 165.100 128.590 165.630 128.615 ;
        RECT 165.100 128.445 165.715 128.590 ;
        RECT 165.470 128.420 165.715 128.445 ;
        RECT 163.435 127.750 165.275 127.775 ;
        RECT 147.215 127.360 153.325 127.530 ;
        RECT 153.760 127.295 156.140 127.625 ;
        RECT 164.010 127.605 165.275 127.750 ;
        RECT 146.775 126.945 148.275 127.115 ;
        RECT 145.720 126.775 146.335 126.945 ;
        RECT 146.165 126.710 146.335 126.775 ;
        RECT 148.105 126.900 148.275 126.945 ;
        RECT 148.105 126.730 153.325 126.900 ;
        RECT 146.165 126.540 147.815 126.710 ;
        RECT 147.645 126.470 147.815 126.540 ;
        RECT 147.645 126.300 148.290 126.470 ;
        RECT 144.905 126.080 145.075 126.185 ;
        RECT 148.120 126.270 148.290 126.300 ;
        RECT 148.120 126.100 153.325 126.270 ;
        RECT 144.905 125.910 147.710 126.080 ;
        RECT 141.725 124.680 142.725 125.680 ;
        RECT 147.540 125.640 147.710 125.910 ;
        RECT 143.965 125.430 147.350 125.600 ;
        RECT 147.540 125.470 153.325 125.640 ;
        RECT 143.965 125.365 144.135 125.430 ;
        RECT 143.605 125.195 144.135 125.365 ;
        RECT 144.760 124.905 146.625 125.075 ;
        RECT 140.405 124.465 140.935 124.550 ;
        RECT 140.405 124.295 141.195 124.465 ;
        RECT 141.025 123.895 141.195 124.295 ;
        RECT 142.375 124.355 142.545 124.680 ;
        RECT 144.760 124.355 144.930 124.905 ;
        RECT 142.375 124.185 144.930 124.355 ;
        RECT 146.455 124.380 146.625 124.905 ;
        RECT 147.180 125.010 147.350 125.430 ;
        RECT 147.180 124.840 153.325 125.010 ;
        RECT 146.455 124.210 153.325 124.380 ;
        RECT 142.015 123.895 144.290 123.920 ;
        RECT 105.585 123.035 106.115 123.205 ;
        RECT 115.820 123.160 116.350 123.330 ;
        RECT 96.600 122.685 97.130 122.855 ;
        RECT 95.965 121.755 96.295 122.180 ;
        RECT 96.775 122.100 96.945 122.685 ;
        RECT 105.770 122.190 105.940 123.035 ;
        RECT 116.005 122.315 116.175 123.160 ;
        RECT 96.730 121.930 101.480 122.100 ;
        RECT 105.745 122.020 110.495 122.190 ;
        RECT 94.610 120.755 96.295 121.755 ;
        RECT 95.965 117.570 96.295 120.755 ;
        RECT 102.140 119.585 102.670 120.115 ;
        RECT 110.930 119.960 111.260 122.270 ;
        RECT 115.895 122.145 120.645 122.315 ;
        RECT 114.740 121.575 115.270 122.105 ;
        RECT 121.080 120.110 121.410 122.395 ;
        RECT 129.160 122.360 129.860 123.800 ;
        RECT 141.025 123.750 144.290 123.895 ;
        RECT 141.025 123.725 142.185 123.750 ;
        RECT 144.120 123.580 153.325 123.750 ;
        RECT 138.510 123.120 139.510 123.520 ;
        RECT 138.510 122.950 153.325 123.120 ;
        RECT 138.510 122.520 139.510 122.950 ;
        RECT 148.575 122.460 153.325 122.490 ;
        RECT 125.130 122.190 129.880 122.360 ;
        RECT 121.080 120.055 122.515 120.110 ;
        RECT 110.930 119.895 112.395 119.960 ;
        RECT 110.930 119.725 112.590 119.895 ;
        RECT 121.080 119.885 122.615 120.055 ;
        RECT 121.080 119.780 122.515 119.885 ;
        RECT 123.900 119.840 124.430 120.370 ;
        RECT 110.930 119.630 112.395 119.725 ;
        RECT 104.580 117.825 105.110 118.355 ;
        RECT 96.730 117.650 101.480 117.820 ;
        RECT 105.745 117.740 110.495 117.910 ;
        RECT 96.800 117.110 96.970 117.650 ;
        RECT 105.785 117.285 105.955 117.740 ;
        RECT 110.930 117.660 111.260 119.630 ;
        RECT 115.895 117.865 120.645 118.035 ;
        RECT 116.280 117.400 116.450 117.865 ;
        RECT 121.080 117.785 121.410 119.780 ;
        RECT 125.130 117.910 129.880 118.080 ;
        RECT 125.135 117.550 125.305 117.910 ;
        RECT 96.340 116.110 97.340 117.110 ;
        RECT 105.325 116.285 106.325 117.285 ;
        RECT 115.820 116.400 116.820 117.400 ;
        RECT 124.865 116.550 125.865 117.550 ;
        RECT 130.315 116.675 130.645 122.440 ;
        RECT 147.035 122.320 153.325 122.460 ;
        RECT 147.035 122.290 148.790 122.320 ;
        RECT 147.035 122.190 147.205 122.290 ;
        RECT 140.405 122.020 147.205 122.190 ;
        RECT 147.600 121.860 148.740 121.875 ;
        RECT 147.600 121.705 153.325 121.860 ;
        RECT 147.600 121.655 147.770 121.705 ;
        RECT 148.575 121.690 153.325 121.705 ;
        RECT 141.460 121.485 147.770 121.655 ;
        RECT 141.460 121.140 141.630 121.485 ;
        RECT 148.575 121.210 153.325 121.230 ;
        RECT 148.060 121.170 153.325 121.210 ;
        RECT 141.045 120.140 142.045 121.140 ;
        RECT 143.185 121.060 153.325 121.170 ;
        RECT 143.185 121.040 148.730 121.060 ;
        RECT 143.185 121.000 148.230 121.040 ;
        RECT 143.185 120.725 143.355 121.000 ;
        RECT 142.740 120.555 143.355 120.725 ;
        RECT 143.840 120.430 153.325 120.600 ;
        RECT 143.840 119.715 144.010 120.430 ;
        RECT 145.305 119.800 153.325 119.970 ;
        RECT 143.120 118.715 144.120 119.715 ;
        RECT 145.305 119.205 145.475 119.800 ;
        RECT 144.845 119.035 145.475 119.205 ;
        RECT 145.025 118.995 145.475 119.035 ;
        RECT 146.015 119.170 153.325 119.340 ;
        RECT 146.015 118.300 146.185 119.170 ;
        RECT 143.995 118.130 146.185 118.300 ;
        RECT 146.625 118.540 153.325 118.710 ;
        RECT 143.995 117.770 144.165 118.130 ;
        RECT 143.120 117.185 144.165 117.770 ;
        RECT 146.625 117.450 146.795 118.540 ;
        RECT 145.230 117.380 146.795 117.450 ;
        RECT 145.050 117.280 146.795 117.380 ;
        RECT 147.245 117.910 153.325 118.080 ;
        RECT 145.050 117.210 145.580 117.280 ;
        RECT 143.120 116.770 144.120 117.185 ;
        RECT 147.245 116.895 147.415 117.910 ;
        RECT 129.940 116.510 130.645 116.675 ;
        RECT 146.185 116.725 147.415 116.895 ;
        RECT 147.735 117.280 153.325 117.450 ;
        RECT 129.940 116.505 130.470 116.510 ;
        RECT 146.185 116.230 146.355 116.725 ;
        RECT 145.390 115.230 146.390 116.230 ;
        RECT 147.735 115.955 147.905 117.280 ;
        RECT 148.575 116.650 153.325 116.820 ;
        RECT 148.960 116.230 149.130 116.650 ;
        RECT 153.760 116.570 154.090 127.295 ;
        RECT 155.140 127.065 156.140 127.295 ;
        RECT 162.405 126.185 163.405 127.185 ;
        RECT 165.105 127.115 165.275 127.605 ;
        RECT 165.545 127.530 165.715 128.420 ;
        RECT 166.065 128.150 166.235 129.475 ;
        RECT 167.210 128.790 167.380 129.695 ;
        RECT 166.920 128.620 171.670 128.790 ;
        RECT 166.920 128.150 171.670 128.160 ;
        RECT 166.065 127.990 171.670 128.150 ;
        RECT 166.065 127.980 167.035 127.990 ;
        RECT 165.545 127.360 171.670 127.530 ;
        RECT 165.105 126.945 166.605 127.115 ;
        RECT 164.050 126.775 164.665 126.945 ;
        RECT 164.495 126.710 164.665 126.775 ;
        RECT 166.435 126.900 166.605 126.945 ;
        RECT 166.435 126.730 171.670 126.900 ;
        RECT 164.495 126.540 166.145 126.710 ;
        RECT 165.975 126.470 166.145 126.540 ;
        RECT 165.975 126.300 166.620 126.470 ;
        RECT 163.235 126.080 163.405 126.185 ;
        RECT 166.450 126.270 166.620 126.300 ;
        RECT 166.450 126.100 171.670 126.270 ;
        RECT 163.235 125.910 166.040 126.080 ;
        RECT 160.055 124.680 161.055 125.680 ;
        RECT 165.870 125.640 166.040 125.910 ;
        RECT 162.295 125.430 165.680 125.600 ;
        RECT 165.870 125.470 171.670 125.640 ;
        RECT 162.295 125.365 162.465 125.430 ;
        RECT 161.935 125.195 162.465 125.365 ;
        RECT 163.090 124.905 164.955 125.075 ;
        RECT 158.735 124.465 159.265 124.550 ;
        RECT 158.735 124.295 159.525 124.465 ;
        RECT 159.355 123.895 159.525 124.295 ;
        RECT 160.705 124.355 160.875 124.680 ;
        RECT 163.090 124.355 163.260 124.905 ;
        RECT 160.705 124.185 163.260 124.355 ;
        RECT 164.785 124.380 164.955 124.905 ;
        RECT 165.510 125.010 165.680 125.430 ;
        RECT 165.510 124.840 171.670 125.010 ;
        RECT 164.785 124.210 171.670 124.380 ;
        RECT 160.345 123.895 162.620 123.920 ;
        RECT 159.355 123.750 162.620 123.895 ;
        RECT 159.355 123.725 160.515 123.750 ;
        RECT 162.450 123.580 171.670 123.750 ;
        RECT 156.840 123.120 157.840 123.540 ;
        RECT 172.105 123.495 172.435 128.870 ;
        RECT 156.840 122.950 171.670 123.120 ;
        RECT 156.840 122.540 157.840 122.950 ;
        RECT 172.105 122.795 173.550 123.495 ;
        RECT 166.920 122.460 171.670 122.490 ;
        RECT 165.365 122.320 171.670 122.460 ;
        RECT 165.365 122.290 167.120 122.320 ;
        RECT 165.365 122.190 165.535 122.290 ;
        RECT 158.735 122.020 165.535 122.190 ;
        RECT 165.930 121.860 167.070 121.875 ;
        RECT 165.930 121.705 171.670 121.860 ;
        RECT 165.930 121.655 166.100 121.705 ;
        RECT 166.920 121.690 171.670 121.705 ;
        RECT 159.790 121.485 166.100 121.655 ;
        RECT 159.790 121.140 159.960 121.485 ;
        RECT 166.920 121.210 171.670 121.230 ;
        RECT 166.390 121.170 171.670 121.210 ;
        RECT 159.375 120.140 160.375 121.140 ;
        RECT 161.515 121.060 171.670 121.170 ;
        RECT 161.515 121.040 167.060 121.060 ;
        RECT 161.515 121.000 166.560 121.040 ;
        RECT 161.515 120.725 161.685 121.000 ;
        RECT 161.070 120.555 161.685 120.725 ;
        RECT 162.170 120.430 171.670 120.600 ;
        RECT 162.170 119.715 162.340 120.430 ;
        RECT 163.635 119.800 171.670 119.970 ;
        RECT 161.450 118.715 162.450 119.715 ;
        RECT 163.635 119.205 163.805 119.800 ;
        RECT 163.175 119.035 163.805 119.205 ;
        RECT 163.355 118.995 163.805 119.035 ;
        RECT 164.345 119.170 171.670 119.340 ;
        RECT 164.345 118.300 164.515 119.170 ;
        RECT 162.325 118.130 164.515 118.300 ;
        RECT 164.955 118.540 171.670 118.710 ;
        RECT 162.325 117.770 162.495 118.130 ;
        RECT 161.450 117.185 162.495 117.770 ;
        RECT 164.955 117.450 165.125 118.540 ;
        RECT 163.560 117.380 165.125 117.450 ;
        RECT 163.380 117.280 165.125 117.380 ;
        RECT 165.575 117.910 171.670 118.080 ;
        RECT 163.380 117.210 163.910 117.280 ;
        RECT 161.450 116.770 162.450 117.185 ;
        RECT 165.575 116.895 165.745 117.910 ;
        RECT 164.515 116.725 165.745 116.895 ;
        RECT 166.065 117.280 171.670 117.450 ;
        RECT 164.515 116.230 164.685 116.725 ;
        RECT 147.310 115.920 147.905 115.955 ;
        RECT 147.130 115.785 147.905 115.920 ;
        RECT 147.130 115.750 147.660 115.785 ;
        RECT 148.545 115.230 149.545 116.230 ;
        RECT 163.720 115.230 164.720 116.230 ;
        RECT 166.065 115.955 166.235 117.280 ;
        RECT 166.920 116.650 171.670 116.820 ;
        RECT 167.290 116.230 167.460 116.650 ;
        RECT 172.105 116.570 172.435 122.795 ;
        RECT 165.640 115.920 166.235 115.955 ;
        RECT 165.460 115.785 166.235 115.920 ;
        RECT 165.460 115.750 165.990 115.785 ;
        RECT 166.875 115.230 167.875 116.230 ;
        RECT 96.600 113.610 97.130 113.780 ;
        RECT 95.965 111.185 96.295 113.115 ;
        RECT 96.775 113.035 96.945 113.610 ;
        RECT 105.585 113.600 106.115 113.770 ;
        RECT 115.820 113.645 116.350 113.815 ;
        RECT 96.730 112.865 101.480 113.035 ;
        RECT 105.760 112.990 105.930 113.600 ;
        RECT 104.580 112.405 105.110 112.935 ;
        RECT 105.745 112.820 110.495 112.990 ;
        RECT 94.240 110.185 96.295 111.185 ;
        RECT 110.930 111.010 111.260 113.070 ;
        RECT 115.995 112.895 116.165 113.645 ;
        RECT 129.410 113.500 129.940 113.505 ;
        RECT 129.230 113.335 129.940 113.500 ;
        RECT 114.740 112.310 115.270 112.840 ;
        RECT 115.895 112.725 120.645 112.895 ;
        RECT 110.930 110.960 112.360 111.010 ;
        RECT 102.160 110.385 102.690 110.915 ;
        RECT 110.930 110.790 112.590 110.960 ;
        RECT 110.930 110.680 112.360 110.790 ;
        RECT 121.080 110.780 121.410 112.975 ;
        RECT 129.230 112.800 129.930 113.335 ;
        RECT 125.175 112.630 129.930 112.800 ;
        RECT 129.230 112.615 129.930 112.630 ;
        RECT 121.080 110.730 122.290 110.780 ;
        RECT 95.965 108.505 96.295 110.185 ;
        RECT 96.730 108.585 101.480 108.755 ;
        RECT 96.800 108.105 96.970 108.585 ;
        RECT 105.745 108.540 110.495 108.710 ;
        RECT 96.340 107.105 97.340 108.105 ;
        RECT 105.785 108.080 105.955 108.540 ;
        RECT 110.930 108.460 111.260 110.680 ;
        RECT 121.080 110.560 122.615 110.730 ;
        RECT 121.080 110.450 122.290 110.560 ;
        RECT 115.895 108.445 120.645 108.615 ;
        RECT 116.280 108.225 116.450 108.445 ;
        RECT 121.080 108.365 121.410 110.450 ;
        RECT 123.920 110.140 124.450 110.670 ;
        RECT 125.185 108.520 125.355 108.540 ;
        RECT 125.175 108.350 129.925 108.520 ;
        RECT 105.325 107.080 106.325 108.080 ;
        RECT 115.820 107.225 116.820 108.225 ;
        RECT 125.185 107.925 125.355 108.350 ;
        RECT 124.460 106.925 125.460 107.925 ;
        RECT 130.360 107.235 130.690 112.880 ;
        RECT 143.495 111.155 144.025 111.685 ;
        RECT 146.770 111.185 147.770 112.185 ;
        RECT 148.410 111.405 148.940 111.575 ;
        RECT 144.815 109.485 145.815 110.460 ;
        RECT 146.480 110.300 147.010 110.325 ;
        RECT 146.480 110.155 147.095 110.300 ;
        RECT 146.850 110.130 147.095 110.155 ;
        RECT 144.815 109.460 146.655 109.485 ;
        RECT 145.390 109.315 146.655 109.460 ;
        RECT 143.785 107.895 144.785 108.895 ;
        RECT 146.485 108.825 146.655 109.315 ;
        RECT 146.925 109.240 147.095 110.130 ;
        RECT 147.445 109.860 147.615 111.185 ;
        RECT 148.590 110.500 148.760 111.405 ;
        RECT 162.145 110.780 162.675 111.310 ;
        RECT 165.370 110.940 166.370 111.940 ;
        RECT 167.060 111.160 167.590 111.330 ;
        RECT 148.270 110.330 153.020 110.500 ;
        RECT 148.270 109.860 153.020 109.870 ;
        RECT 147.445 109.700 153.020 109.860 ;
        RECT 147.445 109.690 148.415 109.700 ;
        RECT 146.925 109.070 153.020 109.240 ;
        RECT 146.485 108.655 147.985 108.825 ;
        RECT 145.430 108.485 146.045 108.655 ;
        RECT 145.875 108.420 146.045 108.485 ;
        RECT 147.815 108.610 147.985 108.655 ;
        RECT 147.815 108.440 153.020 108.610 ;
        RECT 145.875 108.250 147.525 108.420 ;
        RECT 147.355 108.180 147.525 108.250 ;
        RECT 147.355 108.010 148.000 108.180 ;
        RECT 144.615 107.790 144.785 107.895 ;
        RECT 147.830 107.980 148.000 108.010 ;
        RECT 147.830 107.810 153.020 107.980 ;
        RECT 144.615 107.620 147.420 107.790 ;
        RECT 130.070 106.905 130.690 107.235 ;
        RECT 141.435 106.390 142.435 107.390 ;
        RECT 147.250 107.350 147.420 107.620 ;
        RECT 143.675 107.140 147.060 107.310 ;
        RECT 147.250 107.180 153.020 107.350 ;
        RECT 143.675 107.075 143.845 107.140 ;
        RECT 143.315 106.905 143.845 107.075 ;
        RECT 144.470 106.615 146.335 106.785 ;
        RECT 140.115 106.175 140.645 106.260 ;
        RECT 140.115 106.005 140.905 106.175 ;
        RECT 101.650 105.775 102.715 105.870 ;
        RECT 101.650 105.605 102.815 105.775 ;
        RECT 140.735 105.605 140.905 106.005 ;
        RECT 142.085 106.065 142.255 106.390 ;
        RECT 144.470 106.065 144.640 106.615 ;
        RECT 142.085 105.895 144.640 106.065 ;
        RECT 146.165 106.090 146.335 106.615 ;
        RECT 146.890 106.720 147.060 107.140 ;
        RECT 146.890 106.550 153.020 106.720 ;
        RECT 146.165 105.920 153.020 106.090 ;
        RECT 141.725 105.605 144.000 105.630 ;
        RECT 101.650 105.540 102.715 105.605 ;
        RECT 101.650 101.290 101.980 105.540 ;
        RECT 102.415 104.820 102.585 105.540 ;
        RECT 140.735 105.460 144.000 105.605 ;
        RECT 140.735 105.435 141.895 105.460 ;
        RECT 143.830 105.290 153.020 105.460 ;
        RECT 138.220 104.830 139.220 105.250 ;
        RECT 102.405 104.650 108.175 104.820 ;
        RECT 138.220 104.660 153.020 104.830 ;
        RECT 138.220 104.250 139.220 104.660 ;
        RECT 148.270 104.170 153.020 104.200 ;
        RECT 146.745 104.030 153.020 104.170 ;
        RECT 146.745 104.000 148.500 104.030 ;
        RECT 146.745 103.900 146.915 104.000 ;
        RECT 140.115 103.730 146.915 103.900 ;
        RECT 147.310 103.570 148.450 103.585 ;
        RECT 126.205 103.275 126.735 103.450 ;
        RECT 147.310 103.415 153.020 103.570 ;
        RECT 147.310 103.365 147.480 103.415 ;
        RECT 148.270 103.400 153.020 103.415 ;
        RECT 126.205 103.105 134.215 103.275 ;
        RECT 126.205 102.920 126.735 103.105 ;
        RECT 114.460 102.805 115.190 102.810 ;
        RECT 114.280 102.795 115.190 102.805 ;
        RECT 108.815 102.130 109.345 102.660 ;
        RECT 114.280 102.640 121.860 102.795 ;
        RECT 114.280 102.635 114.810 102.640 ;
        RECT 115.070 102.625 121.860 102.640 ;
        RECT 112.130 101.715 121.860 101.885 ;
        RECT 102.405 101.520 108.175 101.540 ;
        RECT 102.395 101.370 108.175 101.520 ;
        RECT 102.395 100.905 102.565 101.370 ;
        RECT 101.935 99.905 102.935 100.905 ;
        RECT 112.130 100.065 112.300 101.715 ;
        RECT 114.460 100.985 115.320 100.990 ;
        RECT 114.280 100.975 115.320 100.985 ;
        RECT 114.280 100.820 121.860 100.975 ;
        RECT 114.280 100.815 114.810 100.820 ;
        RECT 115.070 100.805 121.860 100.820 ;
        RECT 112.130 99.895 121.860 100.065 ;
        RECT 101.650 99.235 102.715 99.265 ;
        RECT 101.650 99.065 102.815 99.235 ;
        RECT 101.650 98.935 102.715 99.065 ;
        RECT 101.650 94.600 101.980 98.935 ;
        RECT 102.405 98.130 102.575 98.935 ;
        RECT 112.130 98.245 112.300 99.895 ;
        RECT 114.460 99.165 115.300 99.170 ;
        RECT 114.280 99.155 115.300 99.165 ;
        RECT 114.280 99.000 121.860 99.155 ;
        RECT 114.280 98.995 114.810 99.000 ;
        RECT 115.070 98.985 121.860 99.000 ;
        RECT 102.405 97.960 108.175 98.130 ;
        RECT 112.130 98.075 121.860 98.245 ;
        RECT 108.835 96.795 109.365 97.325 ;
        RECT 112.130 96.425 112.300 98.075 ;
        RECT 114.290 97.335 115.190 97.350 ;
        RECT 114.290 97.180 121.860 97.335 ;
        RECT 115.070 97.165 121.860 97.180 ;
        RECT 112.130 96.255 121.860 96.425 ;
        RECT 102.405 94.830 108.175 94.850 ;
        RECT 102.395 94.680 108.175 94.830 ;
        RECT 102.395 94.215 102.565 94.680 ;
        RECT 112.130 94.605 112.300 96.255 ;
        RECT 114.290 95.515 114.820 95.525 ;
        RECT 114.290 95.355 121.860 95.515 ;
        RECT 114.470 95.345 121.860 95.355 ;
        RECT 112.130 94.435 121.860 94.605 ;
        RECT 101.935 93.215 102.935 94.215 ;
        RECT 112.130 92.785 112.300 94.435 ;
        RECT 114.470 93.700 115.335 93.710 ;
        RECT 114.290 93.695 115.335 93.700 ;
        RECT 114.290 93.540 121.860 93.695 ;
        RECT 114.290 93.530 114.820 93.540 ;
        RECT 115.070 93.525 121.860 93.540 ;
        RECT 112.130 92.615 121.860 92.785 ;
        RECT 101.650 92.540 102.715 92.610 ;
        RECT 101.650 92.370 102.815 92.540 ;
        RECT 101.650 92.280 102.715 92.370 ;
        RECT 101.650 87.910 101.980 92.280 ;
        RECT 102.410 91.440 102.580 92.280 ;
        RECT 112.130 91.775 112.300 92.615 ;
        RECT 114.280 91.875 115.325 91.890 ;
        RECT 112.700 91.775 112.970 91.860 ;
        RECT 112.130 91.605 112.970 91.775 ;
        RECT 114.280 91.720 121.860 91.875 ;
        RECT 115.070 91.705 121.860 91.720 ;
        RECT 102.405 91.270 108.175 91.440 ;
        RECT 112.130 90.965 112.300 91.605 ;
        RECT 112.700 91.530 112.970 91.605 ;
        RECT 112.130 90.795 121.860 90.965 ;
        RECT 112.130 90.065 112.300 90.795 ;
        RECT 114.555 90.070 114.750 90.185 ;
        RECT 114.555 90.065 115.285 90.070 ;
        RECT 111.985 89.895 112.515 90.065 ;
        RECT 114.290 90.055 115.285 90.065 ;
        RECT 114.290 89.900 121.860 90.055 ;
        RECT 122.275 90.040 122.605 102.875 ;
        RECT 125.005 101.825 134.215 101.995 ;
        RECT 125.055 99.435 125.225 101.825 ;
        RECT 126.205 100.715 126.735 100.935 ;
        RECT 126.205 100.545 134.215 100.715 ;
        RECT 126.205 100.405 126.735 100.545 ;
        RECT 125.055 99.265 134.215 99.435 ;
        RECT 125.055 96.875 125.225 99.265 ;
        RECT 126.205 98.155 126.735 98.330 ;
        RECT 126.205 97.985 134.215 98.155 ;
        RECT 126.205 97.800 126.735 97.985 ;
        RECT 125.055 96.705 134.215 96.875 ;
        RECT 125.055 94.315 125.225 96.705 ;
        RECT 126.205 95.595 126.735 95.800 ;
        RECT 126.205 95.425 134.215 95.595 ;
        RECT 126.205 95.270 126.735 95.425 ;
        RECT 125.055 94.145 134.215 94.315 ;
        RECT 125.055 91.755 125.225 94.145 ;
        RECT 126.205 93.035 126.735 93.155 ;
        RECT 126.205 92.865 134.215 93.035 ;
        RECT 126.205 92.625 126.735 92.865 ;
        RECT 125.055 91.585 134.215 91.755 ;
        RECT 125.055 91.175 125.225 91.585 ;
        RECT 125.055 91.025 125.330 91.175 ;
        RECT 125.060 90.845 125.330 91.025 ;
        RECT 114.290 89.895 114.820 89.900 ;
        RECT 115.070 89.885 121.860 89.900 ;
        RECT 122.255 89.805 122.605 90.040 ;
        RECT 125.085 90.010 125.255 90.845 ;
        RECT 126.205 90.475 126.735 90.680 ;
        RECT 126.205 90.305 134.215 90.475 ;
        RECT 126.205 90.150 126.735 90.305 ;
        RECT 134.630 90.225 134.960 103.355 ;
        RECT 141.170 103.195 147.480 103.365 ;
        RECT 141.170 102.850 141.340 103.195 ;
        RECT 148.270 102.920 153.020 102.940 ;
        RECT 147.770 102.880 153.020 102.920 ;
        RECT 140.755 101.850 141.755 102.850 ;
        RECT 142.895 102.770 153.020 102.880 ;
        RECT 142.895 102.750 148.440 102.770 ;
        RECT 142.895 102.710 147.940 102.750 ;
        RECT 142.895 102.435 143.065 102.710 ;
        RECT 142.450 102.265 143.065 102.435 ;
        RECT 143.550 102.140 153.020 102.310 ;
        RECT 143.550 101.425 143.720 102.140 ;
        RECT 145.015 101.510 153.020 101.680 ;
        RECT 142.830 100.425 143.830 101.425 ;
        RECT 145.015 100.915 145.185 101.510 ;
        RECT 144.555 100.745 145.185 100.915 ;
        RECT 144.735 100.705 145.185 100.745 ;
        RECT 145.725 100.880 153.020 101.050 ;
        RECT 145.725 100.010 145.895 100.880 ;
        RECT 143.705 99.840 145.895 100.010 ;
        RECT 146.335 100.250 153.020 100.420 ;
        RECT 143.705 99.480 143.875 99.840 ;
        RECT 142.830 98.895 143.875 99.480 ;
        RECT 146.335 99.160 146.505 100.250 ;
        RECT 144.940 99.090 146.505 99.160 ;
        RECT 144.760 98.990 146.505 99.090 ;
        RECT 146.955 99.620 153.020 99.790 ;
        RECT 144.760 98.920 145.290 98.990 ;
        RECT 142.830 98.480 143.830 98.895 ;
        RECT 146.955 98.605 147.125 99.620 ;
        RECT 153.455 99.335 153.785 110.580 ;
        RECT 163.465 109.240 164.465 110.215 ;
        RECT 165.130 110.055 165.660 110.080 ;
        RECT 165.130 109.910 165.745 110.055 ;
        RECT 165.500 109.885 165.745 109.910 ;
        RECT 163.465 109.215 165.305 109.240 ;
        RECT 164.040 109.070 165.305 109.215 ;
        RECT 162.435 107.650 163.435 108.650 ;
        RECT 165.135 108.580 165.305 109.070 ;
        RECT 165.575 108.995 165.745 109.885 ;
        RECT 166.095 109.615 166.265 110.940 ;
        RECT 167.240 110.255 167.410 111.160 ;
        RECT 166.925 110.085 171.675 110.255 ;
        RECT 166.925 109.615 171.675 109.625 ;
        RECT 166.095 109.455 171.675 109.615 ;
        RECT 166.095 109.445 167.065 109.455 ;
        RECT 165.575 108.825 171.675 108.995 ;
        RECT 165.135 108.410 166.635 108.580 ;
        RECT 164.080 108.240 164.695 108.410 ;
        RECT 164.525 108.175 164.695 108.240 ;
        RECT 166.465 108.365 166.635 108.410 ;
        RECT 166.465 108.195 171.675 108.365 ;
        RECT 164.525 108.005 166.175 108.175 ;
        RECT 166.005 107.935 166.175 108.005 ;
        RECT 166.005 107.765 166.650 107.935 ;
        RECT 163.265 107.545 163.435 107.650 ;
        RECT 166.480 107.735 166.650 107.765 ;
        RECT 166.480 107.565 171.675 107.735 ;
        RECT 163.265 107.375 166.070 107.545 ;
        RECT 160.085 106.145 161.085 107.145 ;
        RECT 165.900 107.105 166.070 107.375 ;
        RECT 162.325 106.895 165.710 107.065 ;
        RECT 165.900 106.935 171.675 107.105 ;
        RECT 162.325 106.830 162.495 106.895 ;
        RECT 161.965 106.660 162.495 106.830 ;
        RECT 163.120 106.370 164.985 106.540 ;
        RECT 158.765 105.930 159.295 106.015 ;
        RECT 158.765 105.760 159.555 105.930 ;
        RECT 159.385 105.360 159.555 105.760 ;
        RECT 160.735 105.820 160.905 106.145 ;
        RECT 163.120 105.820 163.290 106.370 ;
        RECT 160.735 105.650 163.290 105.820 ;
        RECT 164.815 105.845 164.985 106.370 ;
        RECT 165.540 106.475 165.710 106.895 ;
        RECT 165.540 106.305 171.675 106.475 ;
        RECT 164.815 105.675 171.675 105.845 ;
        RECT 160.375 105.360 162.650 105.385 ;
        RECT 159.385 105.215 162.650 105.360 ;
        RECT 159.385 105.190 160.545 105.215 ;
        RECT 162.480 105.045 171.675 105.215 ;
        RECT 156.870 104.585 157.870 105.020 ;
        RECT 172.110 104.890 172.440 110.335 ;
        RECT 156.870 104.415 171.675 104.585 ;
        RECT 156.870 104.020 157.870 104.415 ;
        RECT 172.110 104.190 173.275 104.890 ;
        RECT 166.925 103.925 171.675 103.955 ;
        RECT 165.395 103.785 171.675 103.925 ;
        RECT 165.395 103.755 167.150 103.785 ;
        RECT 165.395 103.655 165.565 103.755 ;
        RECT 158.765 103.485 165.565 103.655 ;
        RECT 165.960 103.325 167.100 103.340 ;
        RECT 165.960 103.170 171.675 103.325 ;
        RECT 165.960 103.120 166.130 103.170 ;
        RECT 166.925 103.155 171.675 103.170 ;
        RECT 159.820 102.950 166.130 103.120 ;
        RECT 159.820 102.605 159.990 102.950 ;
        RECT 166.925 102.675 171.675 102.695 ;
        RECT 166.420 102.635 171.675 102.675 ;
        RECT 159.405 101.605 160.405 102.605 ;
        RECT 161.545 102.525 171.675 102.635 ;
        RECT 161.545 102.505 167.090 102.525 ;
        RECT 161.545 102.465 166.590 102.505 ;
        RECT 161.545 102.190 161.715 102.465 ;
        RECT 161.100 102.020 161.715 102.190 ;
        RECT 162.200 101.895 171.675 102.065 ;
        RECT 162.200 101.180 162.370 101.895 ;
        RECT 163.665 101.265 171.675 101.435 ;
        RECT 161.480 100.180 162.480 101.180 ;
        RECT 163.665 100.670 163.835 101.265 ;
        RECT 163.205 100.500 163.835 100.670 ;
        RECT 163.385 100.460 163.835 100.500 ;
        RECT 164.375 100.635 171.675 100.805 ;
        RECT 164.375 99.765 164.545 100.635 ;
        RECT 162.355 99.595 164.545 99.765 ;
        RECT 164.985 100.005 171.675 100.175 ;
        RECT 154.645 99.335 155.175 99.450 ;
        RECT 145.895 98.435 147.125 98.605 ;
        RECT 147.445 98.990 153.020 99.160 ;
        RECT 153.455 99.035 155.175 99.335 ;
        RECT 162.355 99.235 162.525 99.595 ;
        RECT 145.895 97.940 146.065 98.435 ;
        RECT 145.100 96.940 146.100 97.940 ;
        RECT 147.445 97.665 147.615 98.990 ;
        RECT 148.270 98.360 153.020 98.530 ;
        RECT 148.670 97.940 148.840 98.360 ;
        RECT 153.455 98.280 153.785 99.035 ;
        RECT 154.645 98.920 155.175 99.035 ;
        RECT 161.480 98.650 162.525 99.235 ;
        RECT 164.985 98.915 165.155 100.005 ;
        RECT 163.590 98.845 165.155 98.915 ;
        RECT 163.410 98.745 165.155 98.845 ;
        RECT 165.605 99.375 171.675 99.545 ;
        RECT 163.410 98.675 163.940 98.745 ;
        RECT 161.480 98.235 162.480 98.650 ;
        RECT 165.605 98.360 165.775 99.375 ;
        RECT 164.545 98.190 165.775 98.360 ;
        RECT 166.095 98.745 171.675 98.915 ;
        RECT 147.020 97.630 147.615 97.665 ;
        RECT 146.840 97.495 147.615 97.630 ;
        RECT 146.840 97.460 147.370 97.495 ;
        RECT 148.255 96.940 149.255 97.940 ;
        RECT 164.545 97.695 164.715 98.190 ;
        RECT 163.750 96.695 164.750 97.695 ;
        RECT 166.095 97.420 166.265 98.745 ;
        RECT 166.925 98.115 171.675 98.285 ;
        RECT 167.320 97.695 167.490 98.115 ;
        RECT 172.110 98.035 172.440 104.190 ;
        RECT 165.670 97.385 166.265 97.420 ;
        RECT 165.490 97.250 166.265 97.385 ;
        RECT 165.490 97.215 166.020 97.250 ;
        RECT 166.905 96.695 167.905 97.695 ;
        RECT 157.755 91.585 158.420 91.755 ;
        RECT 122.255 89.540 122.555 89.805 ;
        RECT 122.255 89.240 122.800 89.540 ;
        RECT 124.880 89.480 125.410 90.010 ;
        RECT 108.815 88.310 109.345 88.840 ;
        RECT 102.395 88.160 102.565 88.165 ;
        RECT 102.395 87.990 108.175 88.160 ;
        RECT 122.500 87.995 122.800 89.240 ;
        RECT 134.635 88.165 134.935 90.225 ;
        RECT 156.855 90.180 157.855 90.650 ;
        RECT 158.250 90.640 158.420 91.585 ;
        RECT 159.105 91.060 160.105 92.060 ;
        RECT 160.760 91.585 161.540 91.755 ;
        RECT 159.840 90.850 160.010 91.060 ;
        RECT 159.840 90.680 161.045 90.850 ;
        RECT 158.250 90.470 159.510 90.640 ;
        RECT 159.340 90.215 159.510 90.470 ;
        RECT 156.855 90.010 158.995 90.180 ;
        RECT 159.340 90.045 160.550 90.215 ;
        RECT 156.855 89.650 157.855 90.010 ;
        RECT 158.825 89.655 158.995 90.010 ;
        RECT 158.825 89.485 160.025 89.655 ;
        RECT 159.855 89.035 160.025 89.485 ;
        RECT 160.380 89.545 160.550 90.045 ;
        RECT 160.875 90.060 161.045 90.680 ;
        RECT 161.370 90.580 161.540 91.585 ;
        RECT 162.105 91.645 163.105 92.060 ;
        RECT 162.105 91.060 163.175 91.645 ;
        RECT 161.370 90.410 162.705 90.580 ;
        RECT 160.875 89.890 162.225 90.060 ;
        RECT 160.380 89.375 161.765 89.545 ;
        RECT 134.635 87.995 134.965 88.165 ;
        RECT 102.395 87.550 102.565 87.990 ;
        RECT 101.935 86.550 102.935 87.550 ;
        RECT 122.385 87.465 122.915 87.995 ;
        RECT 134.540 87.465 135.070 87.995 ;
        RECT 156.520 87.975 157.520 88.975 ;
        RECT 159.855 88.865 161.250 89.035 ;
        RECT 158.310 88.510 159.375 88.680 ;
        RECT 159.205 88.440 159.375 88.510 ;
        RECT 159.205 88.270 160.750 88.440 ;
        RECT 157.190 87.630 157.360 87.975 ;
        RECT 101.650 85.480 102.740 85.810 ;
        RECT 110.565 85.765 111.455 86.655 ;
        RECT 114.695 86.100 115.425 86.105 ;
        RECT 114.515 86.090 115.425 86.100 ;
        RECT 114.515 85.935 122.115 86.090 ;
        RECT 114.515 85.930 115.045 85.935 ;
        RECT 115.325 85.920 122.115 85.935 ;
        RECT 101.650 81.270 101.980 85.480 ;
        RECT 102.210 85.440 102.740 85.480 ;
        RECT 102.405 84.800 102.575 85.440 ;
        RECT 111.950 85.180 112.950 85.660 ;
        RECT 111.950 85.010 122.115 85.180 ;
        RECT 102.405 84.630 108.175 84.800 ;
        RECT 111.950 84.660 112.950 85.010 ;
        RECT 114.695 84.280 115.555 84.285 ;
        RECT 114.515 84.270 115.555 84.280 ;
        RECT 114.515 84.115 122.115 84.270 ;
        RECT 114.515 84.110 115.045 84.115 ;
        RECT 115.325 84.100 122.115 84.115 ;
        RECT 111.950 83.360 112.950 83.775 ;
        RECT 108.835 82.740 109.365 83.270 ;
        RECT 111.950 83.190 122.115 83.360 ;
        RECT 111.950 82.775 112.950 83.190 ;
        RECT 114.695 82.460 115.535 82.465 ;
        RECT 114.515 82.450 115.535 82.460 ;
        RECT 114.515 82.295 122.115 82.450 ;
        RECT 114.515 82.290 115.045 82.295 ;
        RECT 115.325 82.280 122.115 82.295 ;
        RECT 111.950 81.540 112.950 81.950 ;
        RECT 102.395 81.520 102.565 81.540 ;
        RECT 102.395 81.350 108.175 81.520 ;
        RECT 111.950 81.370 122.115 81.540 ;
        RECT 102.395 80.925 102.565 81.350 ;
        RECT 111.950 80.950 112.950 81.370 ;
        RECT 87.805 79.005 89.055 80.255 ;
        RECT 101.935 79.925 102.935 80.925 ;
        RECT 114.525 80.625 115.055 80.640 ;
        RECT 115.325 80.625 122.115 80.630 ;
        RECT 114.525 80.470 122.115 80.625 ;
        RECT 114.705 80.460 122.115 80.470 ;
        RECT 114.705 80.455 115.425 80.460 ;
        RECT 111.950 79.720 112.950 80.075 ;
        RECT 111.950 79.550 122.115 79.720 ;
        RECT 94.375 79.140 94.905 79.310 ;
        RECT 88.180 78.680 88.480 79.005 ;
        RECT 88.180 75.070 88.510 78.680 ;
        RECT 94.550 78.600 94.720 79.140 ;
        RECT 98.950 79.135 99.480 79.305 ;
        RECT 88.985 78.430 94.755 78.600 ;
        RECT 94.550 78.420 94.720 78.430 ;
        RECT 98.305 77.280 98.635 78.680 ;
        RECT 99.125 78.600 99.295 79.135 ;
        RECT 111.950 79.075 112.950 79.550 ;
        RECT 114.525 78.805 115.055 78.820 ;
        RECT 115.325 78.805 122.115 78.810 ;
        RECT 114.525 78.650 122.115 78.805 ;
        RECT 114.705 78.640 122.115 78.650 ;
        RECT 114.705 78.635 115.475 78.640 ;
        RECT 99.110 78.430 104.880 78.600 ;
        RECT 99.125 78.415 99.295 78.430 ;
        RECT 97.550 77.165 98.635 77.280 ;
        RECT 111.950 77.900 112.950 78.255 ;
        RECT 111.950 77.730 122.115 77.900 ;
        RECT 111.950 77.255 112.950 77.730 ;
        RECT 95.535 76.580 96.065 77.110 ;
        RECT 97.450 76.995 98.635 77.165 ;
        RECT 114.705 76.995 115.570 77.005 ;
        RECT 97.550 76.950 98.635 76.995 ;
        RECT 88.985 75.150 94.755 75.320 ;
        RECT 90.320 74.695 90.490 75.150 ;
        RECT 98.305 75.070 98.635 76.950 ;
        RECT 114.525 76.990 115.570 76.995 ;
        RECT 114.525 76.835 122.115 76.990 ;
        RECT 114.525 76.825 115.055 76.835 ;
        RECT 115.325 76.820 122.115 76.835 ;
        RECT 105.595 76.165 106.125 76.695 ;
        RECT 111.950 76.080 112.950 76.515 ;
        RECT 111.950 75.910 122.115 76.080 ;
        RECT 111.950 75.515 112.950 75.910 ;
        RECT 99.110 75.150 104.880 75.320 ;
        RECT 114.515 75.170 115.560 75.185 ;
        RECT 99.130 74.705 99.300 75.150 ;
        RECT 114.515 75.015 122.115 75.170 ;
        RECT 115.325 75.000 122.115 75.015 ;
        RECT 89.860 73.695 90.860 74.695 ;
        RECT 98.670 73.705 99.670 74.705 ;
        RECT 111.950 74.260 112.950 74.680 ;
        RECT 111.950 74.090 122.115 74.260 ;
        RECT 111.950 73.680 112.950 74.090 ;
        RECT 87.805 72.275 89.055 73.525 ;
        RECT 114.790 73.365 114.985 73.480 ;
        RECT 114.790 73.360 115.520 73.365 ;
        RECT 114.525 73.350 115.520 73.360 ;
        RECT 114.525 73.195 122.115 73.350 ;
        RECT 114.525 73.190 115.055 73.195 ;
        RECT 115.325 73.180 122.115 73.195 ;
        RECT 122.530 73.100 122.860 87.465 ;
        RECT 125.205 85.630 125.815 86.300 ;
        RECT 126.205 85.625 126.735 85.805 ;
        RECT 134.635 85.710 134.965 87.465 ;
        RECT 157.190 87.460 160.155 87.630 ;
        RECT 157.450 86.505 159.305 86.510 ;
        RECT 157.270 86.340 159.305 86.505 ;
        RECT 157.270 86.335 157.800 86.340 ;
        RECT 127.445 85.625 134.235 85.630 ;
        RECT 126.205 85.460 134.235 85.625 ;
        RECT 134.635 85.500 134.980 85.710 ;
        RECT 126.205 85.455 127.625 85.460 ;
        RECT 126.205 85.275 126.735 85.455 ;
        RECT 123.485 84.345 124.485 84.775 ;
        RECT 127.445 84.345 134.235 84.350 ;
        RECT 123.485 84.180 134.235 84.345 ;
        RECT 123.485 84.175 127.620 84.180 ;
        RECT 123.485 83.775 124.485 84.175 ;
        RECT 126.130 83.065 126.660 83.240 ;
        RECT 127.445 83.065 134.235 83.070 ;
        RECT 126.130 82.900 134.235 83.065 ;
        RECT 126.130 82.895 127.515 82.900 ;
        RECT 126.130 82.710 126.660 82.895 ;
        RECT 123.425 81.785 124.425 82.205 ;
        RECT 127.445 81.785 134.235 81.790 ;
        RECT 123.425 81.620 134.235 81.785 ;
        RECT 123.425 81.615 127.515 81.620 ;
        RECT 123.425 81.205 124.425 81.615 ;
        RECT 126.125 80.505 126.655 80.685 ;
        RECT 127.445 80.505 134.235 80.510 ;
        RECT 126.125 80.340 134.235 80.505 ;
        RECT 126.125 80.335 127.515 80.340 ;
        RECT 126.125 80.155 126.655 80.335 ;
        RECT 123.535 79.225 124.535 79.700 ;
        RECT 127.445 79.225 134.235 79.230 ;
        RECT 123.535 79.060 134.235 79.225 ;
        RECT 123.535 79.055 127.515 79.060 ;
        RECT 123.535 78.700 124.535 79.055 ;
        RECT 126.165 77.945 126.695 78.120 ;
        RECT 127.445 77.945 134.235 77.950 ;
        RECT 126.165 77.780 134.235 77.945 ;
        RECT 126.165 77.775 127.515 77.780 ;
        RECT 126.165 77.590 126.695 77.775 ;
        RECT 123.535 76.665 124.535 77.090 ;
        RECT 127.445 76.665 134.235 76.670 ;
        RECT 123.535 76.500 134.235 76.665 ;
        RECT 123.535 76.495 127.515 76.500 ;
        RECT 123.535 76.090 124.535 76.495 ;
        RECT 126.140 75.385 126.670 75.560 ;
        RECT 127.445 75.385 134.235 75.390 ;
        RECT 126.140 75.220 134.235 75.385 ;
        RECT 126.140 75.215 127.515 75.220 ;
        RECT 126.140 75.030 126.670 75.215 ;
        RECT 123.535 74.105 124.535 74.605 ;
        RECT 127.445 74.105 134.235 74.110 ;
        RECT 123.535 73.940 134.235 74.105 ;
        RECT 123.535 73.935 127.515 73.940 ;
        RECT 123.535 73.605 124.535 73.935 ;
        RECT 94.395 72.480 94.925 72.650 ;
        RECT 98.950 72.505 99.480 72.675 ;
        RECT 127.445 72.660 134.235 72.830 ;
        RECT 88.185 71.985 88.505 72.275 ;
        RECT 88.180 68.375 88.510 71.985 ;
        RECT 94.570 71.905 94.740 72.480 ;
        RECT 88.985 71.735 94.755 71.905 ;
        RECT 95.505 69.875 96.035 70.405 ;
        RECT 98.305 70.235 98.635 71.985 ;
        RECT 99.125 71.905 99.295 72.505 ;
        RECT 126.615 71.955 127.145 72.135 ;
        RECT 128.205 71.955 128.375 72.660 ;
        RECT 134.650 72.580 134.980 85.500 ;
        RECT 159.135 85.555 159.305 86.340 ;
        RECT 159.985 86.185 160.155 87.460 ;
        RECT 160.580 86.815 160.750 88.270 ;
        RECT 161.080 87.445 161.250 88.865 ;
        RECT 161.595 88.075 161.765 89.375 ;
        RECT 162.055 88.705 162.225 89.890 ;
        RECT 162.535 89.335 162.705 90.410 ;
        RECT 163.005 89.965 163.175 91.060 ;
        RECT 164.645 90.595 165.345 91.755 ;
        RECT 164.090 90.425 170.880 90.595 ;
        RECT 163.005 89.795 170.880 89.965 ;
        RECT 162.535 89.165 170.880 89.335 ;
        RECT 162.055 88.535 170.880 88.705 ;
        RECT 161.595 87.905 170.880 88.075 ;
        RECT 161.080 87.275 170.880 87.445 ;
        RECT 160.580 86.645 170.880 86.815 ;
        RECT 159.985 86.015 170.880 86.185 ;
        RECT 171.295 85.560 171.625 90.675 ;
        RECT 159.135 85.385 170.880 85.555 ;
        RECT 156.520 84.925 157.520 85.355 ;
        RECT 156.520 84.755 170.880 84.925 ;
        RECT 171.295 84.860 173.000 85.560 ;
        RECT 156.520 84.355 157.520 84.755 ;
        RECT 158.975 84.125 170.880 84.295 ;
        RECT 158.975 83.230 159.145 84.125 ;
        RECT 157.450 83.225 159.145 83.230 ;
        RECT 157.270 83.060 159.145 83.225 ;
        RECT 159.865 83.665 164.255 83.675 ;
        RECT 159.865 83.505 170.880 83.665 ;
        RECT 157.270 83.055 157.800 83.060 ;
        RECT 159.865 82.365 160.035 83.505 ;
        RECT 164.090 83.495 170.880 83.505 ;
        RECT 159.070 82.195 160.035 82.365 ;
        RECT 160.475 82.865 170.880 83.035 ;
        RECT 159.070 82.110 159.240 82.195 ;
        RECT 156.935 81.940 159.240 82.110 ;
        RECT 156.935 81.605 157.105 81.940 ;
        RECT 160.475 81.690 160.645 82.865 ;
        RECT 156.520 80.605 157.520 81.605 ;
        RECT 159.680 81.520 160.645 81.690 ;
        RECT 161.000 82.235 170.880 82.405 ;
        RECT 159.680 81.185 159.850 81.520 ;
        RECT 158.310 81.015 159.850 81.185 ;
        RECT 161.000 81.070 161.170 82.235 ;
        RECT 160.220 80.900 161.170 81.070 ;
        RECT 161.585 81.605 170.880 81.775 ;
        RECT 160.220 80.070 160.390 80.900 ;
        RECT 161.585 80.490 161.755 81.605 ;
        RECT 157.195 79.515 158.195 80.000 ;
        RECT 159.230 79.900 160.390 80.070 ;
        RECT 160.760 80.320 161.755 80.490 ;
        RECT 162.075 80.975 170.880 81.145 ;
        RECT 159.230 79.515 159.400 79.900 ;
        RECT 157.195 79.345 159.400 79.515 ;
        RECT 160.760 79.490 160.930 80.320 ;
        RECT 162.075 79.880 162.245 80.975 ;
        RECT 157.195 79.000 158.195 79.345 ;
        RECT 159.895 79.320 160.930 79.490 ;
        RECT 161.280 79.710 162.245 79.880 ;
        RECT 162.635 80.345 170.880 80.515 ;
        RECT 159.895 79.055 160.065 79.320 ;
        RECT 158.805 78.885 160.065 79.055 ;
        RECT 161.280 79.005 161.450 79.710 ;
        RECT 162.635 79.240 162.805 80.345 ;
        RECT 158.805 78.055 158.975 78.885 ;
        RECT 160.445 78.835 161.450 79.005 ;
        RECT 161.790 79.070 162.805 79.240 ;
        RECT 163.295 79.715 170.880 79.885 ;
        RECT 160.445 78.510 160.615 78.835 ;
        RECT 158.310 77.885 158.975 78.055 ;
        RECT 158.490 77.875 158.975 77.885 ;
        RECT 159.605 77.925 160.615 78.510 ;
        RECT 161.790 78.055 161.960 79.070 ;
        RECT 163.295 78.550 163.465 79.715 ;
        RECT 164.090 79.085 170.880 79.255 ;
        RECT 164.900 79.080 165.080 79.085 ;
        RECT 161.390 78.030 161.960 78.055 ;
        RECT 159.605 77.510 160.605 77.925 ;
        RECT 161.210 77.885 161.960 78.030 ;
        RECT 162.335 77.980 163.465 78.550 ;
        RECT 164.910 78.285 165.080 79.080 ;
        RECT 171.295 79.005 171.625 84.860 ;
        RECT 164.730 78.115 165.260 78.285 ;
        RECT 161.210 77.860 161.740 77.885 ;
        RECT 162.335 77.550 163.335 77.980 ;
        RECT 163.320 75.520 163.850 76.050 ;
        RECT 99.110 71.735 104.880 71.905 ;
        RECT 126.615 71.785 128.375 71.955 ;
        RECT 126.615 71.605 127.145 71.785 ;
        RECT 108.410 70.360 108.940 70.690 ;
        RECT 97.550 70.200 98.635 70.235 ;
        RECT 97.450 70.030 98.635 70.200 ;
        RECT 97.550 69.905 98.635 70.030 ;
        RECT 88.985 68.455 94.755 68.625 ;
        RECT 89.970 67.990 90.140 68.455 ;
        RECT 98.305 68.375 98.635 69.905 ;
        RECT 105.615 69.830 106.145 70.360 ;
        RECT 108.610 69.005 108.940 70.360 ;
        RECT 109.510 69.470 110.510 70.470 ;
        RECT 123.405 69.885 124.295 70.775 ;
        RECT 109.210 69.005 109.540 69.050 ;
        RECT 108.610 68.675 109.540 69.005 ;
        RECT 110.010 68.970 110.180 69.470 ;
        RECT 109.955 68.800 116.745 68.970 ;
        RECT 99.110 68.455 104.880 68.625 ;
        RECT 99.115 68.000 99.285 68.455 ;
        RECT 87.805 66.180 89.055 67.430 ;
        RECT 89.510 66.990 90.510 67.990 ;
        RECT 98.655 67.000 99.655 68.000 ;
        RECT 109.210 67.810 109.540 68.675 ;
        RECT 117.115 68.110 117.725 68.780 ;
        RECT 122.660 68.755 122.990 69.225 ;
        RECT 123.840 69.145 124.010 69.885 ;
        RECT 123.405 68.975 130.195 69.145 ;
        RECT 121.590 68.695 122.990 68.755 ;
        RECT 121.490 68.525 122.990 68.695 ;
        RECT 121.590 68.425 122.990 68.525 ;
        RECT 109.955 67.890 116.745 68.060 ;
        RECT 122.660 67.985 122.990 68.425 ;
        RECT 123.405 68.065 130.195 68.235 ;
        RECT 131.165 68.230 131.775 68.900 ;
        RECT 109.970 67.425 110.140 67.890 ;
        RECT 94.355 66.365 94.885 66.535 ;
        RECT 88.190 65.870 88.510 66.180 ;
        RECT 88.180 62.260 88.510 65.870 ;
        RECT 94.530 65.790 94.700 66.365 ;
        RECT 100.140 66.345 100.670 66.515 ;
        RECT 109.510 66.425 110.510 67.425 ;
        RECT 124.050 67.345 124.220 68.065 ;
        RECT 123.870 66.815 124.400 67.345 ;
        RECT 88.985 65.620 94.755 65.790 ;
        RECT 95.505 63.785 96.035 64.315 ;
        RECT 98.305 63.995 98.635 65.870 ;
        RECT 100.315 65.790 100.485 66.345 ;
        RECT 99.110 65.620 104.880 65.790 ;
        RECT 97.450 63.665 98.635 63.995 ;
        RECT 105.615 63.805 106.145 64.335 ;
        RECT 88.985 62.340 94.755 62.510 ;
        RECT 89.970 61.875 90.140 62.340 ;
        RECT 98.305 62.260 98.635 63.665 ;
        RECT 99.150 62.510 99.320 62.520 ;
        RECT 99.110 62.340 104.880 62.510 ;
        RECT 99.150 61.905 99.320 62.340 ;
        RECT 87.975 59.810 89.225 61.060 ;
        RECT 89.510 60.875 90.510 61.875 ;
        RECT 98.690 60.905 99.690 61.905 ;
        RECT 114.070 61.425 114.240 62.095 ;
        RECT 94.395 59.940 94.925 60.110 ;
        RECT 100.140 59.940 100.670 60.110 ;
        RECT 88.195 59.465 88.495 59.810 ;
        RECT 88.180 55.855 88.510 59.465 ;
        RECT 94.570 59.385 94.740 59.940 ;
        RECT 88.985 59.215 94.755 59.385 ;
        RECT 98.305 57.910 98.635 59.465 ;
        RECT 100.315 59.385 100.485 59.940 ;
        RECT 99.110 59.215 104.880 59.385 ;
        RECT 114.070 59.005 114.240 60.885 ;
        RECT 139.135 60.215 139.305 62.095 ;
        RECT 97.550 57.840 98.635 57.910 ;
        RECT 95.505 57.310 96.035 57.840 ;
        RECT 97.450 57.670 98.635 57.840 ;
        RECT 97.550 57.580 98.635 57.670 ;
        RECT 88.985 56.095 94.755 56.105 ;
        RECT 88.980 55.935 94.755 56.095 ;
        RECT 88.980 55.480 89.150 55.935 ;
        RECT 98.305 55.855 98.635 57.580 ;
        RECT 105.615 57.460 106.145 57.990 ;
        RECT 114.070 56.585 114.240 58.465 ;
        RECT 139.135 57.795 139.305 59.675 ;
        RECT 139.135 56.585 139.305 57.255 ;
        RECT 99.105 56.105 99.275 56.115 ;
        RECT 99.105 55.935 104.880 56.105 ;
        RECT 99.105 55.500 99.275 55.935 ;
        RECT 88.520 54.480 89.520 55.480 ;
        RECT 98.645 54.500 99.645 55.500 ;
      LAYER met1 ;
        RECT 138.335 255.745 139.335 255.840 ;
        RECT 61.680 254.745 139.335 255.745 ;
        RECT 61.680 38.025 62.680 254.745 ;
        RECT 113.450 253.945 114.450 254.745 ;
        RECT 138.335 253.945 139.335 254.745 ;
        RECT 90.030 248.305 95.705 253.945 ;
        RECT 108.650 248.445 118.650 253.945 ;
        RECT 136.390 248.535 146.390 253.945 ;
        RECT 148.105 251.655 167.035 252.355 ;
        RECT 90.030 247.605 106.860 248.305 ;
        RECT 90.030 223.850 95.705 247.605 ;
        RECT 104.075 246.285 104.775 247.605 ;
        RECT 104.075 245.585 104.830 246.285 ;
        RECT 104.095 243.240 104.795 245.585 ;
        RECT 111.345 245.380 111.935 246.030 ;
        RECT 105.870 243.660 106.460 244.310 ;
        RECT 104.095 242.540 106.850 243.240 ;
        RECT 104.095 241.385 104.795 242.540 ;
        RECT 104.095 240.685 104.830 241.385 ;
        RECT 111.490 241.375 111.790 245.380 ;
        RECT 115.030 243.890 115.730 248.445 ;
        RECT 116.445 244.590 117.035 245.240 ;
        RECT 143.940 243.890 144.640 248.535 ;
        RECT 145.530 244.590 146.120 245.240 ;
        RECT 114.905 242.880 115.855 243.890 ;
        RECT 143.815 242.880 144.765 243.890 ;
        RECT 111.345 240.725 111.935 241.375 ;
        RECT 116.265 240.785 116.855 241.435 ;
        RECT 145.530 240.805 146.120 241.455 ;
        RECT 104.115 236.810 104.815 240.685 ;
        RECT 105.830 238.850 106.420 239.500 ;
        RECT 104.115 236.110 106.775 236.810 ;
        RECT 104.115 234.150 104.870 236.110 ;
        RECT 111.490 234.980 111.790 240.725 ;
        RECT 148.105 240.495 148.805 251.655 ;
        RECT 151.330 251.065 151.920 251.240 ;
        RECT 146.285 240.480 148.805 240.495 ;
        RECT 116.270 239.675 116.850 240.315 ;
        RECT 117.485 239.795 148.805 240.480 ;
        RECT 149.245 250.765 151.920 251.065 ;
        RECT 149.245 243.870 149.545 250.765 ;
        RECT 151.330 250.590 151.920 250.765 ;
        RECT 156.955 249.785 157.555 251.655 ;
        RECT 159.610 250.985 160.200 251.240 ;
        RECT 156.940 249.135 157.555 249.785 ;
        RECT 149.965 247.970 150.565 248.610 ;
        RECT 155.395 244.800 155.985 245.450 ;
        RECT 151.330 243.870 151.920 244.045 ;
        RECT 149.245 243.570 151.920 243.870 ;
        RECT 117.485 239.780 146.985 239.795 ;
        RECT 117.485 239.710 118.185 239.780 ;
        RECT 111.345 234.330 111.935 234.980 ;
        RECT 104.115 231.885 104.815 234.150 ;
        RECT 105.885 232.905 106.475 233.080 ;
        RECT 111.490 232.905 111.790 234.330 ;
        RECT 105.885 232.605 111.790 232.905 ;
        RECT 105.885 232.430 106.475 232.605 ;
        RECT 104.115 231.185 106.830 231.885 ;
        RECT 104.115 230.160 104.815 231.185 ;
        RECT 104.115 229.460 104.830 230.160 ;
        RECT 111.490 229.935 111.790 232.605 ;
        RECT 111.345 229.285 111.935 229.935 ;
        RECT 105.885 228.085 106.475 228.260 ;
        RECT 111.490 228.085 111.790 229.285 ;
        RECT 105.885 227.785 111.790 228.085 ;
        RECT 105.885 227.610 106.475 227.785 ;
        RECT 106.030 225.330 106.330 227.610 ;
        RECT 105.820 224.690 106.400 225.330 ;
        RECT 90.030 223.800 99.650 223.850 ;
        RECT 90.030 223.150 108.230 223.800 ;
        RECT 90.030 219.120 95.705 223.150 ;
        RECT 96.935 221.890 97.635 223.150 ;
        RECT 98.950 223.100 108.230 223.150 ;
        RECT 106.205 221.015 106.795 221.665 ;
        RECT 105.195 219.665 105.785 219.840 ;
        RECT 106.350 219.665 106.650 221.015 ;
        RECT 106.810 219.665 107.390 219.830 ;
        RECT 105.195 219.365 107.390 219.665 ;
        RECT 105.195 219.190 105.785 219.365 ;
        RECT 90.030 218.420 99.595 219.120 ;
        RECT 90.030 214.545 95.705 218.420 ;
        RECT 96.925 217.435 97.625 218.420 ;
        RECT 106.350 217.210 106.650 219.365 ;
        RECT 106.810 219.190 107.390 219.365 ;
        RECT 106.205 216.560 106.795 217.210 ;
        RECT 105.195 215.150 105.785 215.325 ;
        RECT 106.350 215.150 106.650 216.560 ;
        RECT 105.195 214.850 106.650 215.150 ;
        RECT 105.195 214.675 105.785 214.850 ;
        RECT 90.030 214.530 99.485 214.545 ;
        RECT 90.030 213.880 99.595 214.530 ;
        RECT 90.030 213.845 99.485 213.880 ;
        RECT 90.030 209.005 95.705 213.845 ;
        RECT 96.925 212.835 97.625 213.845 ;
        RECT 106.350 212.515 106.650 214.850 ;
        RECT 107.530 213.435 108.230 223.100 ;
        RECT 108.995 222.005 109.575 222.180 ;
        RECT 116.410 222.005 116.710 239.675 ;
        RECT 135.665 238.180 136.365 239.780 ;
        RECT 133.895 237.480 136.365 238.180 ;
        RECT 128.585 235.385 129.165 236.025 ;
        RECT 128.745 234.995 129.045 235.385 ;
        RECT 128.610 234.345 129.200 234.995 ;
        RECT 128.745 231.925 129.045 234.345 ;
        RECT 130.055 231.925 130.645 232.100 ;
        RECT 128.745 231.625 130.645 231.925 ;
        RECT 128.745 227.720 129.045 231.625 ;
        RECT 130.055 231.450 130.645 231.625 ;
        RECT 135.665 231.075 136.365 237.480 ;
        RECT 133.895 230.375 136.365 231.075 ;
        RECT 135.665 229.275 136.365 230.375 ;
        RECT 149.245 236.895 149.545 243.570 ;
        RECT 151.330 243.395 151.920 243.570 ;
        RECT 149.965 240.795 150.565 241.435 ;
        RECT 155.480 237.735 156.070 238.385 ;
        RECT 151.330 236.895 151.920 237.070 ;
        RECT 149.245 236.595 151.920 236.895 ;
        RECT 149.245 229.885 149.545 236.595 ;
        RECT 151.330 236.420 151.920 236.595 ;
        RECT 149.965 233.845 150.565 234.485 ;
        RECT 155.480 230.855 156.070 231.505 ;
        RECT 151.330 229.885 151.920 230.095 ;
        RECT 149.245 229.585 151.920 229.885 ;
        RECT 128.590 227.070 129.180 227.720 ;
        RECT 128.735 225.095 129.035 227.070 ;
        RECT 148.195 226.770 148.795 227.410 ;
        RECT 130.055 225.095 130.645 225.235 ;
        RECT 128.735 224.795 130.645 225.095 ;
        RECT 128.735 223.980 129.035 224.795 ;
        RECT 130.055 224.585 130.645 224.795 ;
        RECT 148.345 223.980 148.645 226.770 ;
        RECT 128.735 223.680 148.645 223.980 ;
        RECT 128.735 223.675 129.035 223.680 ;
        RECT 149.245 223.000 149.545 229.585 ;
        RECT 151.330 229.445 151.920 229.585 ;
        RECT 156.955 227.605 157.555 249.135 ;
        RECT 157.825 250.845 160.200 250.985 ;
        RECT 157.825 243.790 157.965 250.845 ;
        RECT 159.610 250.590 160.200 250.845 ;
        RECT 166.335 249.660 167.035 251.655 ;
        RECT 165.040 248.960 167.035 249.660 ;
        RECT 158.160 248.110 158.760 248.750 ;
        RECT 159.315 244.800 159.905 245.450 ;
        RECT 159.610 243.790 160.200 244.045 ;
        RECT 157.825 243.650 160.200 243.790 ;
        RECT 157.825 236.885 157.965 243.650 ;
        RECT 159.610 243.395 160.200 243.650 ;
        RECT 166.335 242.895 167.035 248.960 ;
        RECT 165.040 242.195 167.035 242.895 ;
        RECT 158.160 241.030 158.760 241.670 ;
        RECT 159.400 237.735 159.990 238.385 ;
        RECT 159.610 236.885 160.200 237.140 ;
        RECT 157.825 236.745 160.200 236.885 ;
        RECT 157.825 229.905 157.965 236.745 ;
        RECT 159.610 236.490 160.200 236.745 ;
        RECT 164.985 235.700 165.685 235.760 ;
        RECT 166.335 235.700 167.035 242.195 ;
        RECT 164.985 235.000 167.035 235.700 ;
        RECT 158.160 234.160 158.760 234.800 ;
        RECT 159.400 230.855 159.990 231.505 ;
        RECT 159.610 229.905 160.200 230.160 ;
        RECT 157.825 229.765 160.200 229.905 ;
        RECT 149.965 226.820 150.565 227.460 ;
        RECT 155.480 223.695 156.070 224.345 ;
        RECT 157.825 223.000 157.965 229.765 ;
        RECT 159.610 229.510 160.200 229.765 ;
        RECT 166.335 228.280 167.035 235.000 ;
        RECT 172.525 228.280 177.030 253.945 ;
        RECT 165.040 227.580 177.030 228.280 ;
        RECT 158.160 226.820 158.760 227.460 ;
        RECT 159.400 223.695 159.990 224.345 ;
        RECT 149.245 222.700 172.105 223.000 ;
        RECT 108.995 221.705 116.710 222.005 ;
        RECT 108.995 221.540 109.575 221.705 ;
        RECT 110.890 219.070 111.120 220.930 ;
        RECT 171.225 220.730 171.455 220.930 ;
        RECT 171.805 220.730 172.105 222.700 ;
        RECT 171.225 220.590 172.105 220.730 ;
        RECT 171.225 220.280 171.455 220.590 ;
        RECT 110.890 216.650 111.120 218.510 ;
        RECT 171.225 217.860 171.455 219.720 ;
        RECT 110.890 214.230 111.120 216.090 ;
        RECT 171.225 215.440 171.455 217.300 ;
        RECT 172.525 214.880 177.030 227.580 ;
        RECT 171.225 214.230 177.030 214.880 ;
        RECT 107.530 212.735 141.065 213.435 ;
        RECT 106.205 211.865 106.795 212.515 ;
        RECT 105.195 210.545 105.785 210.725 ;
        RECT 106.350 210.545 106.650 211.865 ;
        RECT 105.195 210.245 106.650 210.545 ;
        RECT 105.195 210.075 105.785 210.245 ;
        RECT 90.030 208.960 99.085 209.005 ;
        RECT 90.030 208.310 99.510 208.960 ;
        RECT 90.030 208.305 99.085 208.310 ;
        RECT 90.030 204.525 95.705 208.305 ;
        RECT 96.925 207.290 97.625 208.305 ;
        RECT 106.350 206.805 106.650 210.245 ;
        RECT 140.365 209.580 141.065 212.735 ;
        RECT 157.255 211.235 166.110 211.935 ;
        RECT 141.595 210.575 142.185 211.225 ;
        RECT 140.240 208.570 141.190 209.580 ;
        RECT 157.255 209.310 157.955 211.235 ;
        RECT 159.430 211.065 160.020 211.235 ;
        RECT 143.535 208.610 157.955 209.310 ;
        RECT 165.410 209.975 166.110 211.235 ;
        RECT 172.525 209.975 177.030 214.230 ;
        RECT 165.410 209.275 177.030 209.975 ;
        RECT 106.180 206.155 106.770 206.805 ;
        RECT 90.030 203.825 99.565 204.525 ;
        RECT 104.960 204.475 105.550 205.125 ;
        RECT 90.030 199.870 95.705 203.825 ;
        RECT 97.005 202.675 97.705 203.825 ;
        RECT 106.350 202.495 106.650 206.155 ;
        RECT 106.210 201.845 106.800 202.495 ;
        RECT 98.865 199.870 99.565 199.935 ;
        RECT 90.030 199.170 99.565 199.870 ;
        RECT 104.895 199.840 105.485 200.490 ;
        RECT 73.760 183.690 76.000 183.755 ;
        RECT 90.030 183.690 95.705 199.170 ;
        RECT 96.925 198.185 97.625 199.170 ;
        RECT 106.350 197.895 106.650 201.845 ;
        RECT 140.365 199.620 141.065 208.570 ;
        RECT 141.620 206.605 142.210 207.255 ;
        RECT 141.610 200.515 142.200 201.165 ;
        RECT 140.330 198.610 141.280 199.620 ;
        RECT 144.645 199.390 145.345 208.610 ;
        RECT 158.130 207.755 158.730 208.395 ;
        RECT 159.650 205.800 160.240 205.890 ;
        RECT 157.530 205.500 160.240 205.800 ;
        RECT 146.335 200.980 146.925 201.195 ;
        RECT 157.530 200.980 157.830 205.500 ;
        RECT 159.650 205.240 160.240 205.500 ;
        RECT 159.375 204.490 160.075 204.545 ;
        RECT 159.375 203.790 166.100 204.490 ;
        RECT 165.400 203.420 166.100 203.790 ;
        RECT 172.525 203.420 177.030 209.275 ;
        RECT 165.400 202.745 177.030 203.420 ;
        RECT 165.455 202.720 177.030 202.745 ;
        RECT 146.335 200.680 157.830 200.980 ;
        RECT 158.130 200.965 158.730 201.605 ;
        RECT 146.335 200.545 146.925 200.680 ;
        RECT 143.545 198.690 145.345 199.390 ;
        RECT 157.530 198.585 157.830 200.680 ;
        RECT 159.650 198.585 160.240 198.760 ;
        RECT 157.530 198.285 160.240 198.585 ;
        RECT 159.650 198.110 160.240 198.285 ;
        RECT 106.190 197.245 106.780 197.895 ;
        RECT 138.480 197.105 139.095 197.110 ;
        RECT 138.445 195.740 139.095 197.105 ;
        RECT 141.620 196.615 142.210 197.265 ;
        RECT 104.900 195.090 105.490 195.740 ;
        RECT 107.840 195.040 165.985 195.740 ;
        RECT 138.445 195.030 139.095 195.040 ;
        RECT 165.285 193.270 165.985 195.040 ;
        RECT 98.250 191.410 98.480 193.270 ;
        RECT 163.255 192.620 165.985 193.270 ;
        RECT 98.250 188.990 98.480 190.850 ;
        RECT 163.255 190.200 163.485 192.060 ;
        RECT 98.250 186.570 98.480 188.430 ;
        RECT 163.255 187.780 163.485 189.640 ;
        RECT 98.250 184.150 98.480 186.010 ;
        RECT 163.255 185.360 163.485 187.220 ;
        RECT 73.760 181.690 95.705 183.690 ;
        RECT 98.250 181.730 98.480 183.590 ;
        RECT 163.255 182.940 163.485 184.800 ;
        RECT 73.760 181.555 76.000 181.690 ;
        RECT 90.030 173.910 95.705 181.690 ;
        RECT 98.250 179.310 98.480 181.170 ;
        RECT 163.255 180.520 163.485 182.380 ;
        RECT 165.285 180.845 165.985 192.620 ;
        RECT 172.525 182.690 177.030 202.720 ;
        RECT 190.610 182.690 192.850 182.770 ;
        RECT 98.250 176.890 98.480 178.750 ;
        RECT 163.255 178.100 163.485 179.960 ;
        RECT 98.250 174.470 98.480 176.330 ;
        RECT 163.255 175.680 163.485 177.540 ;
        RECT 163.255 174.470 164.555 175.120 ;
        RECT 163.905 173.910 164.555 174.470 ;
        RECT 90.030 173.260 164.555 173.910 ;
        RECT 90.030 172.945 95.705 173.260 ;
        RECT 165.030 172.945 170.030 180.845 ;
        RECT 172.525 180.690 192.850 182.690 ;
        RECT 172.525 172.945 177.030 180.690 ;
        RECT 190.610 180.570 192.850 180.690 ;
        RECT 167.020 150.420 168.020 172.945 ;
        RECT 66.490 149.420 168.020 150.420 ;
        RECT 66.490 39.500 67.490 149.420 ;
        RECT 81.150 123.195 87.260 145.410 ;
        RECT 96.415 143.160 97.315 143.320 ;
        RECT 105.400 143.170 106.300 143.330 ;
        RECT 115.635 143.170 116.535 143.330 ;
        RECT 96.395 142.520 97.335 143.160 ;
        RECT 105.380 142.530 106.320 143.170 ;
        RECT 115.615 142.530 116.555 143.170 ;
        RECT 124.040 143.145 124.620 143.785 ;
        RECT 129.140 143.695 130.040 143.855 ;
        RECT 96.415 142.360 97.315 142.520 ;
        RECT 105.400 142.370 106.300 142.530 ;
        RECT 115.635 142.370 116.535 142.530 ;
        RECT 94.660 140.645 95.560 140.805 ;
        RECT 94.640 140.005 95.580 140.645 ;
        RECT 111.875 140.500 112.775 140.660 ;
        RECT 121.900 140.500 122.800 140.660 ;
        RECT 94.660 139.845 95.560 140.005 ;
        RECT 102.110 139.710 102.700 140.360 ;
        RECT 111.855 139.860 112.795 140.500 ;
        RECT 121.880 139.860 122.820 140.500 ;
        RECT 124.150 140.155 124.290 143.145 ;
        RECT 129.120 143.055 130.060 143.695 ;
        RECT 129.140 142.895 130.040 143.055 ;
        RECT 132.325 141.580 132.905 141.765 ;
        RECT 176.525 141.580 181.405 145.410 ;
        RECT 132.280 140.880 181.405 141.580 ;
        RECT 96.340 136.175 97.340 137.175 ;
        RECT 96.415 134.310 97.315 134.470 ;
        RECT 96.395 133.670 97.335 134.310 ;
        RECT 96.415 133.510 97.315 133.670 ;
        RECT 102.350 131.485 102.490 139.710 ;
        RECT 111.875 139.700 112.775 139.860 ;
        RECT 121.900 139.700 122.800 139.860 ;
        RECT 123.910 139.505 124.500 140.155 ;
        RECT 132.730 139.875 133.310 140.070 ;
        RECT 132.730 139.735 133.680 139.875 ;
        RECT 104.550 137.745 105.140 138.395 ;
        RECT 102.335 131.285 102.490 131.485 ;
        RECT 94.660 130.850 95.560 131.010 ;
        RECT 94.640 130.210 95.580 130.850 ;
        RECT 102.335 130.250 102.475 131.285 ;
        RECT 94.660 130.050 95.560 130.210 ;
        RECT 102.130 129.600 102.720 130.250 ;
        RECT 96.340 126.265 97.340 127.265 ;
        RECT 87.740 123.195 88.320 123.445 ;
        RECT 81.150 123.055 88.320 123.195 ;
        RECT 96.415 123.090 97.315 123.250 ;
        RECT 81.150 92.200 87.260 123.055 ;
        RECT 87.740 122.805 88.320 123.055 ;
        RECT 96.395 122.450 97.335 123.090 ;
        RECT 96.415 122.290 97.315 122.450 ;
        RECT 94.660 121.490 95.560 121.650 ;
        RECT 94.640 120.850 95.580 121.490 ;
        RECT 94.660 120.690 95.560 120.850 ;
        RECT 102.335 120.175 102.475 129.600 ;
        RECT 104.775 128.465 104.915 137.745 ;
        RECT 114.710 137.715 115.300 138.365 ;
        RECT 105.325 136.210 106.325 137.210 ;
        RECT 114.930 134.035 115.070 137.715 ;
        RECT 115.820 136.150 116.820 137.150 ;
        RECT 124.150 136.820 124.290 139.505 ;
        RECT 132.730 139.430 133.310 139.735 ;
        RECT 133.540 138.930 133.680 139.735 ;
        RECT 133.485 138.280 133.715 138.930 ;
        RECT 124.760 136.820 125.710 137.190 ;
        RECT 124.150 136.680 125.710 136.820 ;
        RECT 129.790 136.785 130.690 136.945 ;
        RECT 124.150 134.035 124.290 136.680 ;
        RECT 124.760 136.180 125.710 136.680 ;
        RECT 129.770 136.145 130.710 136.785 ;
        RECT 129.790 135.985 130.690 136.145 ;
        RECT 133.485 135.860 133.715 137.720 ;
        RECT 174.320 137.070 174.550 138.930 ;
        RECT 114.930 133.895 124.290 134.035 ;
        RECT 105.400 133.210 106.300 133.370 ;
        RECT 105.380 132.570 106.320 133.210 ;
        RECT 105.400 132.410 106.300 132.570 ;
        RECT 114.930 132.170 115.070 133.895 ;
        RECT 115.635 133.230 116.535 133.390 ;
        RECT 115.615 132.590 116.555 133.230 ;
        RECT 115.635 132.430 116.535 132.590 ;
        RECT 114.710 131.520 115.300 132.170 ;
        RECT 111.875 130.150 112.775 130.310 ;
        RECT 111.855 129.510 112.795 130.150 ;
        RECT 111.875 129.350 112.775 129.510 ;
        RECT 104.550 127.815 105.140 128.465 ;
        RECT 102.110 119.525 102.700 120.175 ;
        RECT 96.340 116.110 97.340 117.110 ;
        RECT 96.415 114.015 97.315 114.175 ;
        RECT 96.395 113.375 97.335 114.015 ;
        RECT 96.415 113.215 97.315 113.375 ;
        RECT 94.055 111.005 94.955 111.165 ;
        RECT 94.035 110.365 94.975 111.005 ;
        RECT 102.335 110.975 102.475 119.525 ;
        RECT 104.775 118.415 104.915 127.815 ;
        RECT 105.325 126.300 106.325 127.300 ;
        RECT 105.400 123.440 106.300 123.600 ;
        RECT 105.380 122.800 106.320 123.440 ;
        RECT 105.400 122.640 106.300 122.800 ;
        RECT 114.930 122.165 115.070 131.520 ;
        RECT 121.900 130.150 122.800 130.310 ;
        RECT 124.150 130.190 124.290 133.895 ;
        RECT 129.065 133.695 129.965 133.855 ;
        RECT 129.045 133.055 129.985 133.695 ;
        RECT 133.485 133.440 133.715 135.300 ;
        RECT 174.320 134.650 174.550 136.510 ;
        RECT 176.525 134.095 181.405 140.880 ;
        RECT 174.445 134.090 181.405 134.095 ;
        RECT 174.320 133.440 181.405 134.090 ;
        RECT 174.445 133.395 181.405 133.440 ;
        RECT 129.065 132.895 129.965 133.055 ;
        RECT 176.525 132.895 181.405 133.395 ;
        RECT 172.565 132.195 181.405 132.895 ;
        RECT 143.890 131.720 163.200 131.860 ;
        RECT 121.880 129.510 122.820 130.150 ;
        RECT 123.930 129.540 124.520 130.190 ;
        RECT 143.890 130.130 144.030 131.720 ;
        RECT 163.060 130.725 163.200 131.720 ;
        RECT 143.775 129.860 144.365 130.130 ;
        RECT 136.610 129.720 144.365 129.860 ;
        RECT 121.900 129.350 122.800 129.510 ;
        RECT 115.820 126.255 116.820 127.255 ;
        RECT 124.150 126.810 124.290 129.540 ;
        RECT 124.760 126.810 125.710 127.290 ;
        RECT 129.790 127.265 130.690 127.425 ;
        RECT 124.150 126.670 125.710 126.810 ;
        RECT 115.635 123.565 116.535 123.725 ;
        RECT 115.615 122.925 116.555 123.565 ;
        RECT 115.635 122.765 116.535 122.925 ;
        RECT 114.710 121.515 115.300 122.165 ;
        RECT 111.875 120.130 112.775 120.290 ;
        RECT 111.855 119.490 112.795 120.130 ;
        RECT 111.875 119.330 112.775 119.490 ;
        RECT 104.550 117.765 105.140 118.415 ;
        RECT 104.765 114.825 104.905 117.765 ;
        RECT 105.325 116.285 106.325 117.285 ;
        RECT 114.935 114.825 115.075 121.515 ;
        RECT 121.900 120.290 122.800 120.450 ;
        RECT 124.150 120.430 124.290 126.670 ;
        RECT 124.760 126.280 125.710 126.670 ;
        RECT 129.770 126.625 130.710 127.265 ;
        RECT 129.790 126.465 130.690 126.625 ;
        RECT 129.065 123.865 129.965 124.025 ;
        RECT 129.045 123.225 129.985 123.865 ;
        RECT 129.065 123.065 129.965 123.225 ;
        RECT 121.880 119.650 122.820 120.290 ;
        RECT 123.870 119.780 124.460 120.430 ;
        RECT 121.900 119.490 122.800 119.650 ;
        RECT 124.150 118.525 124.290 119.780 ;
        RECT 124.135 118.385 124.290 118.525 ;
        RECT 115.820 116.400 116.820 117.400 ;
        RECT 104.765 114.685 115.075 114.825 ;
        RECT 104.765 112.995 104.905 114.685 ;
        RECT 105.400 114.005 106.300 114.165 ;
        RECT 105.380 113.365 106.320 114.005 ;
        RECT 105.400 113.205 106.300 113.365 ;
        RECT 104.550 112.345 105.140 112.995 ;
        RECT 114.935 112.900 115.075 114.685 ;
        RECT 115.635 114.050 116.535 114.210 ;
        RECT 115.615 113.410 116.555 114.050 ;
        RECT 115.635 113.250 116.535 113.410 ;
        RECT 114.710 112.250 115.300 112.900 ;
        RECT 111.875 111.195 112.775 111.355 ;
        RECT 102.130 110.710 102.720 110.975 ;
        RECT 102.905 110.710 103.485 110.960 ;
        RECT 102.130 110.570 103.485 110.710 ;
        RECT 94.055 110.205 94.955 110.365 ;
        RECT 102.130 110.325 102.720 110.570 ;
        RECT 102.905 110.320 103.485 110.570 ;
        RECT 111.855 110.555 112.795 111.195 ;
        RECT 121.900 110.965 122.800 111.125 ;
        RECT 111.875 110.395 112.775 110.555 ;
        RECT 121.880 110.325 122.820 110.965 ;
        RECT 124.150 110.730 124.290 118.385 ;
        RECT 124.865 116.550 125.865 117.550 ;
        RECT 129.755 116.910 130.655 117.070 ;
        RECT 129.735 116.270 130.675 116.910 ;
        RECT 129.755 116.110 130.655 116.270 ;
        RECT 129.225 113.740 130.125 113.900 ;
        RECT 129.205 113.100 130.145 113.740 ;
        RECT 129.225 112.940 130.125 113.100 ;
        RECT 136.610 111.115 136.750 129.720 ;
        RECT 143.775 129.480 144.365 129.720 ;
        RECT 147.010 129.475 148.010 130.475 ;
        RECT 148.515 130.100 149.415 130.260 ;
        RECT 148.495 129.460 149.435 130.100 ;
        RECT 162.810 130.075 163.400 130.725 ;
        RECT 165.340 129.475 166.340 130.475 ;
        RECT 166.845 130.100 167.745 130.260 ;
        RECT 166.825 129.460 167.765 130.100 ;
        RECT 148.515 129.300 149.415 129.460 ;
        RECT 166.845 129.300 167.745 129.460 ;
        RECT 146.585 128.850 147.485 129.010 ;
        RECT 164.915 128.850 165.815 129.010 ;
        RECT 145.105 127.750 146.105 128.750 ;
        RECT 146.565 128.210 147.505 128.850 ;
        RECT 146.585 128.050 147.485 128.210 ;
        RECT 144.075 126.185 145.075 127.185 ;
        RECT 145.535 127.180 146.435 127.340 ;
        RECT 145.515 126.540 146.455 127.180 ;
        RECT 155.140 127.065 156.140 128.065 ;
        RECT 163.435 127.750 164.435 128.750 ;
        RECT 164.895 128.210 165.835 128.850 ;
        RECT 164.915 128.050 165.815 128.210 ;
        RECT 145.535 126.380 146.435 126.540 ;
        RECT 162.405 126.185 163.405 127.185 ;
        RECT 163.865 127.180 164.765 127.340 ;
        RECT 163.845 126.540 164.785 127.180 ;
        RECT 163.865 126.380 164.765 126.540 ;
        RECT 140.220 124.785 141.120 124.945 ;
        RECT 140.200 124.145 141.140 124.785 ;
        RECT 141.725 124.680 142.725 125.680 ;
        RECT 143.420 125.600 144.320 125.760 ;
        RECT 143.400 124.960 144.340 125.600 ;
        RECT 143.420 124.800 144.320 124.960 ;
        RECT 158.550 124.785 159.450 124.945 ;
        RECT 158.530 124.145 159.470 124.785 ;
        RECT 160.055 124.680 161.055 125.680 ;
        RECT 161.750 125.600 162.650 125.760 ;
        RECT 161.730 124.960 162.670 125.600 ;
        RECT 161.750 124.800 162.650 124.960 ;
        RECT 140.220 123.985 141.120 124.145 ;
        RECT 158.550 123.985 159.450 124.145 ;
        RECT 138.510 122.520 139.510 123.520 ;
        RECT 140.220 122.425 141.120 122.585 ;
        RECT 156.840 122.540 157.840 123.540 ;
        RECT 176.525 123.495 181.405 132.195 ;
        RECT 172.430 122.795 181.405 123.495 ;
        RECT 158.550 122.425 159.450 122.585 ;
        RECT 140.200 121.785 141.140 122.425 ;
        RECT 158.530 121.785 159.470 122.425 ;
        RECT 140.220 121.625 141.120 121.785 ;
        RECT 158.550 121.625 159.450 121.785 ;
        RECT 141.045 120.140 142.045 121.140 ;
        RECT 142.555 120.960 143.455 121.120 ;
        RECT 142.535 120.320 143.475 120.960 ;
        RECT 142.555 120.160 143.455 120.320 ;
        RECT 159.375 120.140 160.375 121.140 ;
        RECT 160.885 120.960 161.785 121.120 ;
        RECT 160.865 120.320 161.805 120.960 ;
        RECT 160.885 120.160 161.785 120.320 ;
        RECT 143.120 118.715 144.120 119.715 ;
        RECT 144.660 119.440 145.560 119.600 ;
        RECT 144.640 118.800 145.580 119.440 ;
        RECT 144.660 118.640 145.560 118.800 ;
        RECT 161.450 118.715 162.450 119.715 ;
        RECT 162.990 119.440 163.890 119.600 ;
        RECT 162.970 118.800 163.910 119.440 ;
        RECT 162.990 118.640 163.890 118.800 ;
        RECT 143.120 116.770 144.120 117.770 ;
        RECT 144.865 117.615 145.765 117.775 ;
        RECT 144.845 116.975 145.785 117.615 ;
        RECT 144.865 116.815 145.765 116.975 ;
        RECT 161.450 116.770 162.450 117.770 ;
        RECT 163.195 117.615 164.095 117.775 ;
        RECT 163.175 116.975 164.115 117.615 ;
        RECT 163.195 116.815 164.095 116.975 ;
        RECT 145.390 115.230 146.390 116.230 ;
        RECT 146.945 116.155 147.845 116.315 ;
        RECT 146.925 115.515 147.865 116.155 ;
        RECT 146.945 115.355 147.845 115.515 ;
        RECT 148.545 115.230 149.545 116.230 ;
        RECT 163.720 115.230 164.720 116.230 ;
        RECT 165.275 116.155 166.175 116.315 ;
        RECT 165.255 115.515 166.195 116.155 ;
        RECT 165.275 115.355 166.175 115.515 ;
        RECT 166.875 115.230 167.875 116.230 ;
        RECT 143.640 112.880 162.480 113.020 ;
        RECT 143.640 111.745 143.780 112.880 ;
        RECT 143.465 111.115 144.055 111.745 ;
        RECT 146.770 111.185 147.770 112.185 ;
        RECT 148.225 111.810 149.125 111.970 ;
        RECT 148.205 111.170 149.145 111.810 ;
        RECT 162.340 111.370 162.480 112.880 ;
        RECT 136.610 111.095 144.055 111.115 ;
        RECT 136.610 110.975 143.780 111.095 ;
        RECT 148.225 111.010 149.125 111.170 ;
        RECT 121.900 110.165 122.800 110.325 ;
        RECT 123.890 110.080 124.480 110.730 ;
        RECT 96.340 107.105 97.340 108.105 ;
        RECT 105.325 107.080 106.325 108.080 ;
        RECT 115.820 107.225 116.820 108.225 ;
        RECT 124.460 106.925 125.460 107.925 ;
        RECT 129.885 107.390 130.785 107.550 ;
        RECT 129.865 106.750 130.805 107.390 ;
        RECT 129.885 106.590 130.785 106.750 ;
        RECT 102.100 106.010 103.000 106.170 ;
        RECT 102.080 105.370 103.020 106.010 ;
        RECT 102.100 105.210 103.000 105.370 ;
        RECT 108.825 103.425 109.405 104.065 ;
        RECT 109.010 102.720 109.150 103.425 ;
        RECT 124.915 103.255 125.495 103.505 ;
        RECT 126.175 103.255 126.765 103.510 ;
        RECT 114.095 103.040 114.995 103.200 ;
        RECT 124.915 103.115 126.765 103.255 ;
        RECT 108.785 102.070 109.375 102.720 ;
        RECT 114.075 102.400 115.015 103.040 ;
        RECT 124.915 102.865 125.495 103.115 ;
        RECT 126.175 102.860 126.765 103.115 ;
        RECT 114.095 102.240 114.995 102.400 ;
        RECT 101.935 99.905 102.935 100.905 ;
        RECT 102.100 99.470 103.000 99.630 ;
        RECT 102.080 98.830 103.020 99.470 ;
        RECT 102.100 98.670 103.000 98.830 ;
        RECT 109.025 97.385 109.165 102.070 ;
        RECT 114.095 101.220 114.995 101.380 ;
        RECT 114.075 100.580 115.015 101.220 ;
        RECT 126.400 100.995 126.540 102.860 ;
        RECT 114.095 100.420 114.995 100.580 ;
        RECT 126.175 100.345 126.765 100.995 ;
        RECT 114.095 99.400 114.995 99.560 ;
        RECT 114.075 98.760 115.015 99.400 ;
        RECT 114.095 98.600 114.995 98.760 ;
        RECT 126.400 98.390 126.540 100.345 ;
        RECT 114.105 97.585 115.005 97.745 ;
        RECT 126.175 97.740 126.765 98.390 ;
        RECT 108.805 96.735 109.395 97.385 ;
        RECT 114.085 96.945 115.025 97.585 ;
        RECT 114.105 96.785 115.005 96.945 ;
        RECT 98.385 93.800 98.965 94.030 ;
        RECT 95.695 93.660 98.965 93.800 ;
        RECT 81.150 92.185 88.255 92.200 ;
        RECT 81.150 91.545 88.545 92.185 ;
        RECT 81.150 91.500 88.255 91.545 ;
        RECT 81.150 81.525 87.260 91.500 ;
        RECT 81.150 80.825 88.545 81.525 ;
        RECT 81.150 79.970 87.260 80.825 ;
        RECT 87.775 79.970 89.085 80.315 ;
        RECT 81.150 79.270 89.085 79.970 ;
        RECT 94.190 79.545 95.090 79.705 ;
        RECT 81.150 73.390 87.260 79.270 ;
        RECT 87.775 78.945 89.085 79.270 ;
        RECT 94.170 78.905 95.110 79.545 ;
        RECT 94.190 78.745 95.090 78.905 ;
        RECT 95.695 77.170 95.835 93.660 ;
        RECT 98.385 93.390 98.965 93.660 ;
        RECT 101.935 93.215 102.935 94.215 ;
        RECT 102.100 92.775 103.000 92.935 ;
        RECT 102.080 92.135 103.020 92.775 ;
        RECT 102.100 91.975 103.000 92.135 ;
        RECT 109.010 88.900 109.150 96.735 ;
        RECT 114.105 95.760 115.005 95.920 ;
        RECT 126.400 95.860 126.540 97.740 ;
        RECT 114.085 95.120 115.025 95.760 ;
        RECT 126.175 95.210 126.765 95.860 ;
        RECT 114.105 94.960 115.005 95.120 ;
        RECT 114.105 93.935 115.005 94.095 ;
        RECT 114.085 93.295 115.025 93.935 ;
        RECT 114.105 93.135 115.005 93.295 ;
        RECT 126.400 93.215 126.540 95.210 ;
        RECT 126.175 92.565 126.765 93.215 ;
        RECT 114.095 92.125 114.995 92.285 ;
        RECT 114.075 91.485 115.015 92.125 ;
        RECT 114.095 91.325 114.995 91.485 ;
        RECT 126.400 90.740 126.540 92.565 ;
        RECT 111.800 90.300 112.700 90.460 ;
        RECT 114.105 90.300 115.005 90.460 ;
        RECT 111.780 89.660 112.720 90.300 ;
        RECT 114.085 89.660 115.025 90.300 ;
        RECT 126.175 90.090 126.765 90.740 ;
        RECT 123.595 89.815 124.175 90.080 ;
        RECT 124.850 89.815 125.440 90.070 ;
        RECT 123.595 89.675 125.440 89.815 ;
        RECT 111.800 89.500 112.700 89.660 ;
        RECT 114.105 89.500 115.005 89.660 ;
        RECT 123.595 89.440 124.175 89.675 ;
        RECT 124.850 89.420 125.440 89.675 ;
        RECT 136.610 89.345 136.750 110.975 ;
        RECT 162.115 110.720 162.705 111.370 ;
        RECT 165.370 110.940 166.370 111.940 ;
        RECT 166.875 111.565 167.775 111.725 ;
        RECT 166.855 110.925 167.795 111.565 ;
        RECT 166.875 110.765 167.775 110.925 ;
        RECT 146.295 110.560 147.195 110.720 ;
        RECT 144.815 109.460 145.815 110.460 ;
        RECT 146.275 109.920 147.215 110.560 ;
        RECT 164.945 110.315 165.845 110.475 ;
        RECT 146.295 109.760 147.195 109.920 ;
        RECT 163.465 109.215 164.465 110.215 ;
        RECT 164.925 109.675 165.865 110.315 ;
        RECT 164.945 109.515 165.845 109.675 ;
        RECT 143.785 107.895 144.785 108.895 ;
        RECT 145.245 108.890 146.145 109.050 ;
        RECT 145.225 108.250 146.165 108.890 ;
        RECT 145.245 108.090 146.145 108.250 ;
        RECT 162.435 107.650 163.435 108.650 ;
        RECT 163.895 108.645 164.795 108.805 ;
        RECT 163.875 108.005 164.815 108.645 ;
        RECT 163.895 107.845 164.795 108.005 ;
        RECT 139.930 106.495 140.830 106.655 ;
        RECT 139.910 105.855 140.850 106.495 ;
        RECT 141.435 106.390 142.435 107.390 ;
        RECT 143.130 107.310 144.030 107.470 ;
        RECT 143.110 106.670 144.050 107.310 ;
        RECT 143.130 106.510 144.030 106.670 ;
        RECT 158.580 106.250 159.480 106.410 ;
        RECT 139.930 105.695 140.830 105.855 ;
        RECT 158.560 105.610 159.500 106.250 ;
        RECT 160.085 106.145 161.085 107.145 ;
        RECT 161.780 107.065 162.680 107.225 ;
        RECT 161.760 106.425 162.700 107.065 ;
        RECT 161.780 106.265 162.680 106.425 ;
        RECT 158.580 105.450 159.480 105.610 ;
        RECT 138.220 104.250 139.220 105.250 ;
        RECT 139.930 104.135 140.830 104.295 ;
        RECT 139.910 103.495 140.850 104.135 ;
        RECT 156.870 104.020 157.870 105.020 ;
        RECT 176.525 104.890 181.405 122.795 ;
        RECT 172.715 104.190 181.405 104.890 ;
        RECT 158.580 103.890 159.480 104.050 ;
        RECT 139.930 103.335 140.830 103.495 ;
        RECT 158.560 103.250 159.500 103.890 ;
        RECT 158.580 103.090 159.480 103.250 ;
        RECT 140.755 101.850 141.755 102.850 ;
        RECT 142.265 102.670 143.165 102.830 ;
        RECT 142.245 102.030 143.185 102.670 ;
        RECT 142.265 101.870 143.165 102.030 ;
        RECT 159.405 101.605 160.405 102.605 ;
        RECT 160.915 102.425 161.815 102.585 ;
        RECT 160.895 101.785 161.835 102.425 ;
        RECT 160.915 101.625 161.815 101.785 ;
        RECT 142.830 100.425 143.830 101.425 ;
        RECT 144.370 101.150 145.270 101.310 ;
        RECT 144.350 100.510 145.290 101.150 ;
        RECT 144.370 100.350 145.270 100.510 ;
        RECT 161.480 100.180 162.480 101.180 ;
        RECT 163.020 100.905 163.920 101.065 ;
        RECT 163.000 100.265 163.940 100.905 ;
        RECT 163.020 100.105 163.920 100.265 ;
        RECT 142.830 98.480 143.830 99.480 ;
        RECT 144.575 99.325 145.475 99.485 ;
        RECT 144.555 98.685 145.495 99.325 ;
        RECT 154.615 99.135 155.205 99.510 ;
        RECT 144.575 98.525 145.475 98.685 ;
        RECT 145.100 96.940 146.100 97.940 ;
        RECT 146.655 97.865 147.555 98.025 ;
        RECT 146.635 97.225 147.575 97.865 ;
        RECT 146.655 97.065 147.555 97.225 ;
        RECT 148.255 96.940 149.255 97.940 ;
        RECT 154.560 95.045 155.260 99.135 ;
        RECT 161.480 98.235 162.480 99.235 ;
        RECT 163.225 99.080 164.125 99.240 ;
        RECT 163.205 98.440 164.145 99.080 ;
        RECT 163.225 98.280 164.125 98.440 ;
        RECT 163.750 96.695 164.750 97.695 ;
        RECT 165.305 97.620 166.205 97.780 ;
        RECT 165.285 96.980 166.225 97.620 ;
        RECT 165.305 96.820 166.205 96.980 ;
        RECT 166.905 96.695 167.905 97.695 ;
        RECT 176.525 95.045 181.405 104.190 ;
        RECT 154.560 94.345 181.405 95.045 ;
        RECT 154.590 93.675 155.290 94.345 ;
        RECT 126.310 89.205 136.750 89.345 ;
        RECT 152.105 92.975 155.290 93.675 ;
        RECT 108.785 88.250 109.375 88.900 ;
        RECT 126.310 88.865 126.450 89.205 ;
        RECT 110.885 88.725 126.450 88.865 ;
        RECT 101.935 86.550 102.935 87.550 ;
        RECT 102.025 85.845 102.925 86.005 ;
        RECT 102.005 85.205 102.945 85.845 ;
        RECT 102.025 85.045 102.925 85.205 ;
        RECT 109.025 83.330 109.165 88.250 ;
        RECT 110.885 86.715 111.025 88.725 ;
        RECT 152.105 88.080 152.805 92.975 ;
        RECT 157.570 91.990 158.470 92.150 ;
        RECT 157.550 91.350 158.490 91.990 ;
        RECT 157.570 91.190 158.470 91.350 ;
        RECT 159.105 91.060 160.105 92.060 ;
        RECT 160.575 91.990 161.475 92.150 ;
        RECT 160.555 91.350 161.495 91.990 ;
        RECT 160.575 91.190 161.475 91.350 ;
        RECT 162.105 91.060 163.105 92.060 ;
        RECT 164.545 91.990 165.445 92.150 ;
        RECT 164.525 91.350 165.465 91.990 ;
        RECT 164.545 91.190 165.445 91.350 ;
        RECT 156.855 89.650 157.855 90.650 ;
        RECT 122.355 87.380 152.805 88.080 ;
        RECT 156.520 87.975 157.520 88.975 ;
        RECT 158.125 88.915 159.025 89.075 ;
        RECT 158.105 88.275 159.045 88.915 ;
        RECT 158.125 88.115 159.025 88.275 ;
        RECT 110.535 85.705 111.485 86.715 ;
        RECT 114.330 86.335 115.230 86.495 ;
        RECT 110.940 84.155 111.080 85.705 ;
        RECT 114.310 85.695 115.250 86.335 ;
        RECT 123.595 86.035 124.175 86.330 ;
        RECT 125.215 86.035 125.805 86.290 ;
        RECT 123.595 85.895 125.805 86.035 ;
        RECT 111.950 84.660 112.950 85.660 ;
        RECT 114.330 85.535 115.230 85.695 ;
        RECT 123.595 85.690 124.175 85.895 ;
        RECT 125.215 85.640 125.805 85.895 ;
        RECT 126.120 85.890 126.820 87.380 ;
        RECT 157.085 86.740 157.985 86.900 ;
        RECT 157.065 86.100 158.005 86.740 ;
        RECT 157.085 85.940 157.985 86.100 ;
        RECT 126.060 85.610 126.820 85.890 ;
        RECT 126.060 85.470 126.935 85.610 ;
        RECT 176.525 85.600 181.405 94.345 ;
        RECT 126.060 85.190 126.820 85.470 ;
        RECT 114.330 84.515 115.230 84.675 ;
        RECT 110.645 83.515 111.225 84.155 ;
        RECT 114.310 83.875 115.250 84.515 ;
        RECT 108.805 82.680 109.395 83.330 ;
        RECT 111.950 82.775 112.950 83.775 ;
        RECT 114.330 83.715 115.230 83.875 ;
        RECT 123.485 83.775 124.485 84.775 ;
        RECT 126.325 83.300 126.465 85.190 ;
        RECT 156.520 84.355 157.520 85.355 ;
        RECT 172.355 84.900 181.405 85.600 ;
        RECT 157.085 83.460 157.985 83.620 ;
        RECT 114.330 82.695 115.230 82.855 ;
        RECT 114.310 82.055 115.250 82.695 ;
        RECT 126.100 82.650 126.690 83.300 ;
        RECT 157.065 82.820 158.005 83.460 ;
        RECT 157.085 82.660 157.985 82.820 ;
        RECT 111.950 80.950 112.950 81.950 ;
        RECT 114.330 81.895 115.230 82.055 ;
        RECT 123.425 81.205 124.425 82.205 ;
        RECT 101.935 79.925 102.935 80.925 ;
        RECT 114.340 80.875 115.240 81.035 ;
        RECT 114.320 80.235 115.260 80.875 ;
        RECT 126.320 80.745 126.460 82.650 ;
        RECT 114.340 80.075 115.240 80.235 ;
        RECT 126.095 80.095 126.685 80.745 ;
        RECT 156.520 80.605 157.520 81.605 ;
        RECT 158.125 81.420 159.025 81.580 ;
        RECT 158.105 80.780 159.045 81.420 ;
        RECT 158.125 80.620 159.025 80.780 ;
        RECT 98.765 79.540 99.665 79.700 ;
        RECT 98.745 78.900 99.685 79.540 ;
        RECT 111.950 79.075 112.950 80.075 ;
        RECT 114.340 79.055 115.240 79.215 ;
        RECT 98.765 78.740 99.665 78.900 ;
        RECT 114.320 78.415 115.260 79.055 ;
        RECT 123.535 78.700 124.535 79.700 ;
        RECT 114.340 78.255 115.240 78.415 ;
        RECT 97.265 77.400 98.165 77.560 ;
        RECT 95.505 76.520 96.095 77.170 ;
        RECT 97.245 76.760 98.185 77.400 ;
        RECT 111.950 77.255 112.950 78.255 ;
        RECT 126.360 78.180 126.500 80.095 ;
        RECT 157.195 79.000 158.195 80.000 ;
        RECT 158.125 78.290 159.025 78.450 ;
        RECT 126.135 77.530 126.725 78.180 ;
        RECT 158.105 77.650 159.045 78.290 ;
        RECT 114.340 77.230 115.240 77.390 ;
        RECT 97.265 76.600 98.165 76.760 ;
        RECT 89.860 73.695 90.860 74.695 ;
        RECT 87.775 73.390 89.085 73.585 ;
        RECT 81.150 72.690 89.085 73.390 ;
        RECT 94.210 72.885 95.110 73.045 ;
        RECT 81.150 66.895 87.260 72.690 ;
        RECT 87.775 72.215 89.085 72.690 ;
        RECT 94.190 72.245 95.130 72.885 ;
        RECT 94.210 72.085 95.110 72.245 ;
        RECT 95.695 71.095 95.835 76.520 ;
        RECT 105.565 76.105 106.155 76.755 ;
        RECT 114.320 76.590 115.260 77.230 ;
        RECT 98.670 73.705 99.670 74.705 ;
        RECT 98.765 72.910 99.665 73.070 ;
        RECT 98.745 72.270 99.685 72.910 ;
        RECT 98.765 72.110 99.665 72.270 ;
        RECT 105.805 71.095 105.945 76.105 ;
        RECT 111.950 75.515 112.950 76.515 ;
        RECT 114.340 76.430 115.240 76.590 ;
        RECT 123.535 76.090 124.535 77.090 ;
        RECT 126.335 75.620 126.475 77.530 ;
        RECT 158.125 77.490 159.025 77.650 ;
        RECT 159.605 77.510 160.605 78.510 ;
        RECT 161.025 78.265 161.925 78.425 ;
        RECT 161.005 77.625 161.945 78.265 ;
        RECT 161.025 77.465 161.925 77.625 ;
        RECT 162.335 77.550 163.335 78.550 ;
        RECT 164.545 78.520 165.445 78.680 ;
        RECT 164.525 77.880 165.465 78.520 ;
        RECT 176.525 78.500 181.405 84.900 ;
        RECT 176.250 78.450 181.405 78.500 ;
        RECT 164.545 77.720 165.445 77.880 ;
        RECT 175.885 77.810 181.405 78.450 ;
        RECT 176.250 77.800 181.405 77.810 ;
        RECT 114.330 75.420 115.230 75.580 ;
        RECT 114.310 74.780 115.250 75.420 ;
        RECT 126.110 74.970 126.700 75.620 ;
        RECT 163.290 75.460 163.880 76.110 ;
        RECT 111.950 73.680 112.950 74.680 ;
        RECT 114.330 74.620 115.230 74.780 ;
        RECT 114.340 73.595 115.240 73.755 ;
        RECT 123.535 73.605 124.535 74.605 ;
        RECT 114.320 72.955 115.260 73.595 ;
        RECT 114.340 72.795 115.240 72.955 ;
        RECT 123.630 72.570 124.210 72.740 ;
        RECT 120.600 72.270 125.225 72.570 ;
        RECT 95.695 70.950 95.840 71.095 ;
        RECT 105.805 70.950 105.950 71.095 ;
        RECT 95.700 70.465 95.840 70.950 ;
        RECT 95.475 69.815 96.065 70.465 ;
        RECT 97.265 70.435 98.165 70.595 ;
        RECT 87.775 66.895 89.085 67.490 ;
        RECT 89.510 66.990 90.510 67.990 ;
        RECT 81.150 66.195 89.085 66.895 ;
        RECT 94.170 66.770 95.070 66.930 ;
        RECT 73.760 64.665 76.000 64.675 ;
        RECT 81.150 64.665 87.260 66.195 ;
        RECT 87.775 66.120 89.085 66.195 ;
        RECT 94.150 66.130 95.090 66.770 ;
        RECT 94.170 65.970 95.070 66.130 ;
        RECT 73.760 62.665 87.260 64.665 ;
        RECT 95.700 64.375 95.840 69.815 ;
        RECT 97.245 69.795 98.185 70.435 ;
        RECT 105.810 70.420 105.950 70.950 ;
        RECT 108.225 70.845 109.125 71.005 ;
        RECT 97.265 69.635 98.165 69.795 ;
        RECT 105.585 69.770 106.175 70.420 ;
        RECT 108.205 70.205 109.145 70.845 ;
        RECT 108.225 70.045 109.125 70.205 ;
        RECT 98.655 67.000 99.655 68.000 ;
        RECT 99.955 66.750 100.855 66.910 ;
        RECT 99.935 66.110 100.875 66.750 ;
        RECT 99.955 65.950 100.855 66.110 ;
        RECT 105.810 64.395 105.950 69.770 ;
        RECT 109.510 69.470 110.510 70.470 ;
        RECT 117.125 68.710 117.715 68.770 ;
        RECT 117.125 68.120 117.855 68.710 ;
        RECT 109.510 66.425 110.510 67.425 ;
        RECT 95.475 63.725 96.065 64.375 ;
        RECT 97.265 64.150 98.165 64.310 ;
        RECT 73.760 62.475 76.000 62.665 ;
        RECT 81.150 60.670 87.260 62.665 ;
        RECT 87.945 60.670 89.255 61.120 ;
        RECT 89.510 60.875 90.510 61.875 ;
        RECT 81.150 59.970 89.255 60.670 ;
        RECT 94.210 60.345 95.110 60.505 ;
        RECT 81.150 52.085 87.260 59.970 ;
        RECT 87.945 59.750 89.255 59.970 ;
        RECT 94.190 59.705 95.130 60.345 ;
        RECT 94.210 59.545 95.110 59.705 ;
        RECT 95.700 57.900 95.840 63.725 ;
        RECT 97.245 63.510 98.185 64.150 ;
        RECT 105.585 63.745 106.175 64.395 ;
        RECT 97.265 63.350 98.165 63.510 ;
        RECT 98.690 60.905 99.690 61.905 ;
        RECT 99.955 60.345 100.855 60.505 ;
        RECT 99.935 59.705 100.875 60.345 ;
        RECT 99.955 59.545 100.855 59.705 ;
        RECT 97.265 58.075 98.165 58.235 ;
        RECT 95.475 57.250 96.065 57.900 ;
        RECT 97.245 57.435 98.185 58.075 ;
        RECT 105.810 58.050 105.950 63.745 ;
        RECT 107.435 61.435 114.270 62.085 ;
        RECT 97.265 57.275 98.165 57.435 ;
        RECT 105.585 57.400 106.175 58.050 ;
        RECT 88.520 54.480 89.520 55.480 ;
        RECT 95.700 53.015 95.840 57.250 ;
        RECT 98.645 54.500 99.645 55.500 ;
        RECT 105.810 53.015 105.950 57.400 ;
        RECT 95.700 52.875 105.950 53.015 ;
        RECT 107.435 52.085 108.085 61.435 ;
        RECT 114.040 59.015 114.270 60.875 ;
        RECT 114.040 56.595 114.270 58.455 ;
        RECT 81.150 51.435 108.085 52.085 ;
        RECT 81.150 45.620 87.260 51.435 ;
        RECT 117.155 50.885 117.855 68.120 ;
        RECT 120.600 67.220 120.900 72.270 ;
        RECT 123.630 72.100 124.210 72.270 ;
        RECT 124.925 71.360 125.225 72.270 ;
        RECT 126.280 71.940 126.420 74.970 ;
        RECT 163.515 74.630 163.655 75.460 ;
        RECT 163.215 73.990 163.795 74.630 ;
        RECT 126.585 71.940 127.175 72.195 ;
        RECT 126.280 71.800 127.175 71.940 ;
        RECT 126.585 71.545 127.175 71.800 ;
        RECT 123.375 69.825 124.325 70.835 ;
        RECT 124.860 70.720 125.440 71.360 ;
        RECT 121.305 68.930 122.205 69.090 ;
        RECT 121.285 68.290 122.225 68.930 ;
        RECT 121.305 68.130 122.205 68.290 ;
        RECT 123.840 67.220 124.430 67.405 ;
        RECT 120.600 66.920 124.430 67.220 ;
        RECT 123.840 66.755 124.430 66.920 ;
        RECT 107.880 45.605 117.880 50.885 ;
        RECT 131.110 50.700 131.810 68.960 ;
        RECT 139.105 60.225 139.335 62.085 ;
        RECT 139.105 57.805 139.335 59.665 ;
        RECT 139.105 56.595 140.315 57.245 ;
        RECT 139.665 53.455 140.315 56.595 ;
        RECT 147.730 53.455 148.730 53.630 ;
        RECT 139.665 52.805 148.730 53.455 ;
        RECT 139.665 50.870 140.315 52.805 ;
        RECT 147.730 52.630 148.730 52.805 ;
        RECT 176.525 51.860 181.405 77.800 ;
        RECT 190.610 51.860 192.850 51.940 ;
        RECT 121.820 45.625 131.820 50.700 ;
        RECT 138.785 45.630 148.785 50.870 ;
        RECT 176.525 49.860 192.850 51.860 ;
        RECT 116.235 41.235 117.235 45.605 ;
        RECT 130.025 43.140 131.025 45.625 ;
        RECT 144.175 45.080 145.175 45.630 ;
        RECT 176.525 45.620 181.405 49.860 ;
        RECT 190.610 49.740 192.850 49.860 ;
        RECT 191.090 45.080 192.370 45.220 ;
        RECT 144.175 44.080 192.370 45.080 ;
        RECT 191.090 43.980 192.370 44.080 ;
        RECT 130.025 43.010 181.470 43.140 ;
        RECT 130.025 42.140 182.040 43.010 ;
        RECT 180.760 41.770 182.040 42.140 ;
        RECT 116.235 41.090 159.225 41.235 ;
        RECT 116.235 40.235 160.105 41.090 ;
        RECT 158.825 39.850 160.105 40.235 ;
        RECT 66.490 39.425 137.460 39.500 ;
        RECT 66.490 38.875 137.765 39.425 ;
        RECT 66.530 38.500 137.765 38.875 ;
        RECT 136.485 38.185 137.765 38.500 ;
        RECT 61.680 37.885 114.725 38.025 ;
        RECT 61.680 37.025 115.590 37.885 ;
        RECT 114.310 36.645 115.590 37.025 ;
      LAYER met2 ;
        RECT 149.900 247.905 150.630 248.675 ;
        RECT 158.095 248.045 158.825 248.815 ;
        RECT 155.400 245.345 155.980 245.445 ;
        RECT 159.320 245.345 159.900 245.445 ;
        RECT 116.450 245.065 117.030 245.235 ;
        RECT 145.535 245.065 146.115 245.235 ;
        RECT 155.400 245.205 159.900 245.345 ;
        RECT 116.450 244.765 147.645 245.065 ;
        RECT 155.400 244.805 155.980 245.205 ;
        RECT 116.450 244.595 117.030 244.765 ;
        RECT 145.535 244.595 146.115 244.765 ;
        RECT 105.875 244.105 106.455 244.305 ;
        RECT 105.875 243.805 113.180 244.105 ;
        RECT 105.875 243.665 106.455 243.805 ;
        RECT 105.835 239.265 106.415 239.495 ;
        RECT 112.880 239.265 113.180 243.805 ;
        RECT 116.270 241.280 116.850 241.430 ;
        RECT 145.535 241.280 146.115 241.450 ;
        RECT 116.270 240.980 146.115 241.280 ;
        RECT 116.270 240.790 116.850 240.980 ;
        RECT 145.535 240.810 146.115 240.980 ;
        RECT 116.410 240.315 116.710 240.790 ;
        RECT 116.270 239.675 116.850 240.315 ;
        RECT 105.835 238.965 128.985 239.265 ;
        RECT 105.835 238.855 106.415 238.965 ;
        RECT 128.685 236.025 128.985 238.965 ;
        RECT 128.585 235.385 129.165 236.025 ;
        RECT 105.545 224.425 106.675 225.595 ;
        RECT 108.995 221.540 109.575 222.180 ;
        RECT 106.810 219.660 107.390 219.830 ;
        RECT 109.140 219.660 109.440 221.540 ;
        RECT 106.810 219.360 109.440 219.660 ;
        RECT 106.810 219.190 107.390 219.360 ;
        RECT 141.600 211.050 142.180 211.220 ;
        RECT 141.600 211.010 145.900 211.050 ;
        RECT 147.345 211.010 147.645 244.765 ;
        RECT 149.900 240.730 150.630 241.500 ;
        RECT 155.485 238.130 156.065 238.380 ;
        RECT 157.630 238.130 157.770 245.205 ;
        RECT 159.320 244.805 159.900 245.205 ;
        RECT 158.095 240.965 158.825 241.735 ;
        RECT 159.405 238.130 159.985 238.380 ;
        RECT 155.485 237.990 159.985 238.130 ;
        RECT 155.485 237.740 156.065 237.990 ;
        RECT 149.900 233.780 150.630 234.550 ;
        RECT 155.485 231.250 156.065 231.500 ;
        RECT 157.630 231.250 157.770 237.990 ;
        RECT 159.405 237.740 159.985 237.990 ;
        RECT 158.095 234.095 158.825 234.865 ;
        RECT 159.405 231.250 159.985 231.500 ;
        RECT 155.485 231.110 159.985 231.250 ;
        RECT 155.485 230.860 156.065 231.110 ;
        RECT 148.130 226.705 148.860 227.475 ;
        RECT 149.900 226.755 150.630 227.525 ;
        RECT 149.900 224.090 150.630 224.495 ;
        RECT 155.485 224.090 156.065 224.340 ;
        RECT 157.630 224.090 157.770 231.110 ;
        RECT 159.405 230.860 159.985 231.110 ;
        RECT 158.095 226.755 158.825 227.525 ;
        RECT 159.405 224.090 159.985 224.340 ;
        RECT 149.900 223.950 159.985 224.090 ;
        RECT 149.900 223.725 150.630 223.950 ;
        RECT 155.485 223.700 156.065 223.950 ;
        RECT 159.405 223.700 159.985 223.950 ;
        RECT 141.600 210.750 147.645 211.010 ;
        RECT 141.600 210.580 142.180 210.750 ;
        RECT 145.600 210.710 147.645 210.750 ;
        RECT 141.625 207.035 142.205 207.250 ;
        RECT 138.585 206.735 142.205 207.035 ;
        RECT 105.110 205.160 105.810 205.165 ;
        RECT 104.880 204.460 107.600 205.160 ;
        RECT 104.900 200.480 105.480 200.485 ;
        RECT 106.900 200.480 107.600 204.460 ;
        RECT 104.900 199.845 107.600 200.480 ;
        RECT 104.940 199.780 107.600 199.845 ;
        RECT 104.905 195.720 105.800 195.735 ;
        RECT 106.900 195.720 107.600 199.780 ;
        RECT 138.585 197.105 138.885 206.735 ;
        RECT 141.625 206.610 142.205 206.735 ;
        RECT 141.615 200.990 142.195 201.160 ;
        RECT 145.600 200.990 145.900 210.710 ;
        RECT 158.065 207.690 158.795 208.460 ;
        RECT 146.340 200.990 146.920 201.190 ;
        RECT 141.615 200.690 146.920 200.990 ;
        RECT 158.065 200.900 158.795 201.670 ;
        RECT 141.615 200.520 142.195 200.690 ;
        RECT 146.340 200.550 146.920 200.690 ;
        RECT 138.480 197.090 139.060 197.105 ;
        RECT 141.625 197.090 142.205 197.260 ;
        RECT 138.480 196.790 142.205 197.090 ;
        RECT 138.480 196.465 139.060 196.790 ;
        RECT 141.625 196.620 142.205 196.790 ;
        RECT 107.780 195.720 108.480 195.735 ;
        RECT 104.845 195.020 108.480 195.720 ;
        RECT 73.695 181.490 76.065 183.820 ;
        RECT 190.545 180.505 192.915 182.835 ;
        RECT 104.520 144.045 133.380 144.185 ;
        RECT 96.415 143.130 97.315 143.320 ;
        RECT 93.960 142.430 97.315 143.130 ;
        RECT 93.960 140.805 94.660 142.430 ;
        RECT 96.415 142.360 97.315 142.430 ;
        RECT 104.520 142.920 104.660 144.045 ;
        RECT 105.400 142.920 106.300 143.330 ;
        RECT 104.520 142.780 106.300 142.920 ;
        RECT 93.960 139.845 95.560 140.805 ;
        RECT 93.960 134.455 94.660 139.845 ;
        RECT 96.275 136.090 97.405 137.260 ;
        RECT 96.415 134.455 97.315 134.470 ;
        RECT 93.960 133.755 97.315 134.455 ;
        RECT 93.960 131.010 94.660 133.755 ;
        RECT 96.285 133.720 97.315 133.755 ;
        RECT 96.415 133.510 97.315 133.720 ;
        RECT 104.520 132.870 104.660 142.780 ;
        RECT 105.400 142.370 106.300 142.780 ;
        RECT 114.705 142.920 114.845 144.045 ;
        RECT 115.635 142.920 116.535 143.330 ;
        RECT 123.965 143.080 124.695 143.850 ;
        RECT 129.140 143.795 130.040 143.855 ;
        RECT 129.140 143.095 132.095 143.795 ;
        RECT 114.705 142.780 116.535 142.920 ;
        RECT 129.140 142.895 130.040 143.095 ;
        RECT 111.875 140.530 112.775 140.660 ;
        RECT 111.855 139.700 112.775 140.530 ;
        RECT 105.260 136.125 106.390 137.295 ;
        RECT 105.400 132.870 106.300 133.370 ;
        RECT 104.510 132.730 106.300 132.870 ;
        RECT 93.960 130.050 95.560 131.010 ;
        RECT 87.740 123.435 88.320 123.445 ;
        RECT 93.960 123.435 94.660 130.050 ;
        RECT 96.275 126.180 97.405 127.350 ;
        RECT 87.740 123.250 96.865 123.435 ;
        RECT 87.740 122.805 97.315 123.250 ;
        RECT 104.520 123.190 104.660 132.730 ;
        RECT 105.400 132.410 106.300 132.730 ;
        RECT 111.855 130.310 112.555 139.700 ;
        RECT 114.705 132.890 114.845 142.780 ;
        RECT 115.635 142.370 116.535 142.780 ;
        RECT 131.395 141.840 132.095 143.095 ;
        RECT 131.395 141.140 132.965 141.840 ;
        RECT 121.900 139.700 122.800 140.660 ;
        RECT 115.755 136.065 116.885 137.235 ;
        RECT 115.635 132.890 116.535 133.390 ;
        RECT 114.705 132.750 116.535 132.890 ;
        RECT 111.855 129.350 112.775 130.310 ;
        RECT 105.260 126.215 106.390 127.385 ;
        RECT 105.400 123.190 106.300 123.600 ;
        RECT 104.510 123.050 106.300 123.190 ;
        RECT 88.030 122.735 97.315 122.805 ;
        RECT 93.960 121.650 94.660 122.735 ;
        RECT 96.415 122.290 97.315 122.735 ;
        RECT 93.960 120.690 95.560 121.650 ;
        RECT 93.960 114.005 94.660 120.690 ;
        RECT 96.275 116.025 97.405 117.195 ;
        RECT 96.415 114.005 97.315 114.175 ;
        RECT 93.960 113.305 97.315 114.005 ;
        RECT 104.520 113.725 104.660 123.050 ;
        RECT 105.400 122.640 106.300 123.050 ;
        RECT 111.855 120.290 112.555 129.350 ;
        RECT 114.705 123.315 114.845 132.750 ;
        RECT 115.635 132.430 116.535 132.750 ;
        RECT 122.000 130.310 122.700 139.700 ;
        RECT 129.790 136.815 130.690 136.945 ;
        RECT 129.775 135.985 130.690 136.815 ;
        RECT 129.775 135.845 130.475 135.985 ;
        RECT 131.395 135.845 132.095 141.140 ;
        RECT 132.265 141.125 132.965 141.140 ;
        RECT 133.240 140.070 133.380 144.045 ;
        RECT 132.730 139.680 133.380 140.070 ;
        RECT 132.730 139.430 133.310 139.680 ;
        RECT 129.135 135.145 132.095 135.845 ;
        RECT 129.135 133.855 129.835 135.145 ;
        RECT 129.065 132.895 129.965 133.855 ;
        RECT 121.900 129.350 122.800 130.310 ;
        RECT 115.755 126.170 116.885 127.340 ;
        RECT 115.635 123.315 116.535 123.725 ;
        RECT 114.705 123.175 116.535 123.315 ;
        RECT 111.855 119.330 112.775 120.290 ;
        RECT 105.260 116.200 106.390 117.370 ;
        RECT 105.400 113.725 106.300 114.165 ;
        RECT 104.520 113.585 106.300 113.725 ;
        RECT 93.960 111.165 94.660 113.305 ;
        RECT 96.415 113.215 97.315 113.305 ;
        RECT 105.400 113.205 106.300 113.585 ;
        RECT 111.855 111.355 112.555 119.330 ;
        RECT 114.705 113.755 114.845 123.175 ;
        RECT 115.635 122.765 116.535 123.175 ;
        RECT 122.000 120.450 122.700 129.350 ;
        RECT 129.790 126.465 130.690 127.425 ;
        RECT 129.890 125.570 130.590 126.465 ;
        RECT 131.395 125.570 132.095 135.145 ;
        RECT 172.500 132.160 173.230 132.930 ;
        RECT 146.490 131.020 167.345 131.160 ;
        RECT 146.490 129.010 146.630 131.020 ;
        RECT 146.945 129.390 148.075 130.560 ;
        RECT 148.835 130.260 148.975 131.020 ;
        RECT 148.515 129.300 149.415 130.260 ;
        RECT 145.040 127.665 146.170 128.835 ;
        RECT 146.490 128.460 147.485 129.010 ;
        RECT 146.585 128.050 147.485 128.460 ;
        RECT 129.110 124.870 132.095 125.570 ;
        RECT 140.600 126.445 143.515 126.585 ;
        RECT 140.600 124.945 140.740 126.445 ;
        RECT 129.110 124.025 129.810 124.870 ;
        RECT 129.065 123.065 129.965 124.025 ;
        RECT 121.900 119.490 122.800 120.450 ;
        RECT 115.755 116.315 116.885 117.485 ;
        RECT 115.635 113.755 116.535 114.210 ;
        RECT 114.705 113.615 116.535 113.755 ;
        RECT 115.635 113.250 116.535 113.615 ;
        RECT 93.960 110.335 94.955 111.165 ;
        RECT 94.055 110.205 94.955 110.335 ;
        RECT 102.830 110.255 103.560 111.025 ;
        RECT 111.855 110.395 112.775 111.355 ;
        RECT 122.000 111.125 122.700 119.490 ;
        RECT 124.800 116.465 125.930 117.635 ;
        RECT 129.755 116.110 130.655 117.070 ;
        RECT 129.930 115.375 130.630 116.110 ;
        RECT 131.395 115.375 132.095 124.870 ;
        RECT 140.220 123.985 141.120 124.945 ;
        RECT 141.660 124.595 142.790 125.765 ;
        RECT 143.375 125.760 143.515 126.445 ;
        RECT 144.010 126.100 145.140 127.270 ;
        RECT 145.535 126.930 146.435 127.340 ;
        RECT 146.875 126.930 147.015 128.050 ;
        RECT 145.535 126.790 147.015 126.930 ;
        RECT 145.535 126.380 146.435 126.790 ;
        RECT 143.375 125.545 144.320 125.760 ;
        RECT 145.915 125.545 146.055 126.380 ;
        RECT 143.375 125.405 146.055 125.545 ;
        RECT 143.375 125.210 144.320 125.405 ;
        RECT 143.420 124.800 144.320 125.210 ;
        RECT 138.445 122.435 139.575 123.605 ;
        RECT 140.600 122.585 140.740 123.985 ;
        RECT 140.220 122.175 141.120 122.585 ;
        RECT 140.180 121.625 141.120 122.175 ;
        RECT 140.180 119.395 140.320 121.625 ;
        RECT 140.980 120.055 142.110 121.225 ;
        RECT 142.555 120.675 143.455 121.120 ;
        RECT 142.555 120.535 145.180 120.675 ;
        RECT 142.555 120.160 143.455 120.535 ;
        RECT 142.700 119.395 142.840 120.160 ;
        RECT 140.180 119.255 142.840 119.395 ;
        RECT 142.195 116.115 142.335 119.255 ;
        RECT 143.055 118.630 144.185 119.800 ;
        RECT 145.040 119.600 145.180 120.535 ;
        RECT 144.660 118.640 145.560 119.600 ;
        RECT 143.055 116.685 144.185 117.855 ;
        RECT 144.865 117.365 145.765 117.775 ;
        RECT 144.780 116.815 145.765 117.365 ;
        RECT 144.780 116.115 144.920 116.815 ;
        RECT 142.195 115.975 144.920 116.115 ;
        RECT 129.295 114.675 132.095 115.375 ;
        RECT 129.295 113.900 129.995 114.675 ;
        RECT 129.225 112.940 130.125 113.900 ;
        RECT 96.275 107.020 97.405 108.190 ;
        RECT 105.260 106.995 106.390 108.165 ;
        RECT 102.100 106.150 103.000 106.170 ;
        RECT 101.370 106.010 103.000 106.150 ;
        RECT 101.370 99.585 101.510 106.010 ;
        RECT 102.100 105.210 103.000 106.010 ;
        RECT 111.855 105.160 112.555 110.395 ;
        RECT 121.900 110.165 122.800 111.125 ;
        RECT 115.755 107.140 116.885 108.310 ;
        RECT 122.000 105.160 122.700 110.165 ;
        RECT 124.395 106.840 125.525 108.010 ;
        RECT 129.885 106.590 130.785 107.550 ;
        RECT 130.050 105.160 130.750 106.590 ;
        RECT 131.395 105.160 132.095 114.675 ;
        RECT 143.845 114.375 143.985 115.975 ;
        RECT 145.325 115.145 146.455 116.315 ;
        RECT 146.945 115.355 147.845 116.315 ;
        RECT 147.325 114.375 147.465 115.355 ;
        RECT 148.480 115.145 149.610 116.315 ;
        RECT 143.845 114.235 147.465 114.375 ;
        RECT 154.590 112.625 154.730 131.020 ;
        RECT 164.820 129.010 164.960 131.020 ;
        RECT 165.275 129.390 166.405 130.560 ;
        RECT 167.205 130.260 167.345 131.020 ;
        RECT 166.845 129.300 167.745 130.260 ;
        RECT 155.075 126.980 156.205 128.150 ;
        RECT 163.370 127.665 164.500 128.835 ;
        RECT 164.820 128.460 165.815 129.010 ;
        RECT 164.915 128.050 165.815 128.460 ;
        RECT 158.930 126.445 161.845 126.585 ;
        RECT 158.930 124.945 159.070 126.445 ;
        RECT 158.550 123.985 159.450 124.945 ;
        RECT 159.990 124.595 161.120 125.765 ;
        RECT 161.705 125.760 161.845 126.445 ;
        RECT 162.340 126.100 163.470 127.270 ;
        RECT 163.865 126.930 164.765 127.340 ;
        RECT 165.205 126.930 165.345 128.050 ;
        RECT 163.865 126.790 165.345 126.930 ;
        RECT 163.865 126.380 164.765 126.790 ;
        RECT 161.705 125.545 162.650 125.760 ;
        RECT 164.245 125.545 164.385 126.380 ;
        RECT 161.705 125.405 164.385 125.545 ;
        RECT 161.705 125.210 162.650 125.405 ;
        RECT 161.750 124.800 162.650 125.210 ;
        RECT 156.775 122.455 157.905 123.625 ;
        RECT 158.930 122.585 159.070 123.985 ;
        RECT 158.550 122.175 159.450 122.585 ;
        RECT 158.510 121.625 159.450 122.175 ;
        RECT 158.510 119.395 158.650 121.625 ;
        RECT 159.310 120.055 160.440 121.225 ;
        RECT 160.885 120.675 161.785 121.120 ;
        RECT 160.885 120.535 163.510 120.675 ;
        RECT 160.885 120.160 161.785 120.535 ;
        RECT 161.030 119.395 161.170 120.160 ;
        RECT 158.510 119.255 161.170 119.395 ;
        RECT 160.525 116.115 160.665 119.255 ;
        RECT 161.385 118.630 162.515 119.800 ;
        RECT 163.370 119.600 163.510 120.535 ;
        RECT 162.990 118.640 163.890 119.600 ;
        RECT 161.385 116.685 162.515 117.855 ;
        RECT 163.195 117.365 164.095 117.775 ;
        RECT 163.110 116.815 164.095 117.365 ;
        RECT 163.110 116.115 163.250 116.815 ;
        RECT 160.525 115.975 163.250 116.115 ;
        RECT 162.175 114.375 162.315 115.975 ;
        RECT 163.655 115.145 164.785 116.315 ;
        RECT 165.275 115.355 166.175 116.315 ;
        RECT 165.655 114.375 165.795 115.355 ;
        RECT 166.810 115.145 167.940 116.315 ;
        RECT 162.175 114.235 165.795 114.375 ;
        RECT 146.415 112.485 167.335 112.625 ;
        RECT 146.415 110.720 146.555 112.485 ;
        RECT 146.705 111.100 147.835 112.270 ;
        RECT 148.430 111.970 148.570 112.485 ;
        RECT 148.225 111.010 149.125 111.970 ;
        RECT 144.750 109.375 145.880 110.545 ;
        RECT 146.295 109.760 147.195 110.720 ;
        RECT 164.850 110.475 164.990 112.485 ;
        RECT 165.305 110.855 166.435 112.025 ;
        RECT 167.195 111.725 167.335 112.485 ;
        RECT 166.875 110.765 167.775 111.725 ;
        RECT 140.310 108.155 143.225 108.295 ;
        RECT 140.310 106.655 140.450 108.155 ;
        RECT 139.930 105.695 140.830 106.655 ;
        RECT 141.370 106.305 142.500 107.475 ;
        RECT 143.085 107.470 143.225 108.155 ;
        RECT 143.720 107.810 144.850 108.980 ;
        RECT 145.245 108.640 146.145 109.050 ;
        RECT 146.585 108.640 146.725 109.760 ;
        RECT 163.400 109.130 164.530 110.300 ;
        RECT 164.850 109.925 165.845 110.475 ;
        RECT 164.945 109.515 165.845 109.925 ;
        RECT 145.245 108.500 146.725 108.640 ;
        RECT 145.245 108.090 146.145 108.500 ;
        RECT 143.085 107.255 144.030 107.470 ;
        RECT 145.625 107.255 145.765 108.090 ;
        RECT 143.085 107.115 145.765 107.255 ;
        RECT 158.960 107.910 161.875 108.050 ;
        RECT 143.085 106.920 144.030 107.115 ;
        RECT 143.130 106.510 144.030 106.920 ;
        RECT 158.960 106.410 159.100 107.910 ;
        RECT 111.855 104.460 132.095 105.160 ;
        RECT 108.750 103.360 109.480 104.130 ;
        RECT 113.480 102.790 113.620 104.460 ;
        RECT 114.095 102.790 114.995 103.200 ;
        RECT 124.855 102.865 125.555 104.460 ;
        RECT 138.155 104.165 139.285 105.335 ;
        RECT 140.310 104.295 140.450 105.695 ;
        RECT 158.580 105.450 159.480 106.410 ;
        RECT 160.020 106.060 161.150 107.230 ;
        RECT 161.735 107.225 161.875 107.910 ;
        RECT 162.370 107.565 163.500 108.735 ;
        RECT 163.895 108.395 164.795 108.805 ;
        RECT 165.235 108.395 165.375 109.515 ;
        RECT 163.895 108.255 165.375 108.395 ;
        RECT 163.895 107.845 164.795 108.255 ;
        RECT 161.735 107.010 162.680 107.225 ;
        RECT 164.275 107.010 164.415 107.845 ;
        RECT 161.735 106.870 164.415 107.010 ;
        RECT 161.735 106.675 162.680 106.870 ;
        RECT 161.780 106.265 162.680 106.675 ;
        RECT 139.930 103.885 140.830 104.295 ;
        RECT 156.805 103.935 157.935 105.105 ;
        RECT 158.960 104.050 159.100 105.450 ;
        RECT 139.890 103.335 140.830 103.885 ;
        RECT 158.580 103.640 159.480 104.050 ;
        RECT 113.480 102.650 114.995 102.790 ;
        RECT 101.870 99.820 103.000 100.990 ;
        RECT 113.480 100.820 113.620 102.650 ;
        RECT 114.095 102.240 114.995 102.650 ;
        RECT 114.095 100.820 114.995 101.380 ;
        RECT 113.480 100.680 114.995 100.820 ;
        RECT 139.890 100.730 140.030 103.335 ;
        RECT 158.540 103.090 159.480 103.640 ;
        RECT 140.690 101.765 141.820 102.935 ;
        RECT 142.265 102.010 143.165 102.830 ;
        RECT 142.265 101.870 144.890 102.010 ;
        RECT 142.410 100.730 142.550 101.870 ;
        RECT 102.100 99.585 103.000 99.630 ;
        RECT 101.370 99.445 103.000 99.585 ;
        RECT 98.310 93.325 99.040 94.095 ;
        RECT 101.370 92.865 101.510 99.445 ;
        RECT 102.100 98.670 103.000 99.445 ;
        RECT 113.480 99.170 113.620 100.680 ;
        RECT 114.095 100.420 114.995 100.680 ;
        RECT 135.815 100.590 142.550 100.730 ;
        RECT 114.095 99.170 114.995 99.560 ;
        RECT 113.480 99.030 114.995 99.170 ;
        RECT 113.480 97.305 113.620 99.030 ;
        RECT 114.095 98.600 114.995 99.030 ;
        RECT 114.105 97.305 115.005 97.745 ;
        RECT 113.480 97.165 115.005 97.305 ;
        RECT 113.480 95.500 113.620 97.165 ;
        RECT 114.105 96.785 115.005 97.165 ;
        RECT 114.105 95.500 115.005 95.920 ;
        RECT 113.480 95.360 115.005 95.500 ;
        RECT 101.870 93.130 103.000 94.300 ;
        RECT 113.480 93.675 113.620 95.360 ;
        RECT 114.105 94.960 115.005 95.360 ;
        RECT 114.105 93.675 115.005 94.095 ;
        RECT 113.480 93.535 115.005 93.675 ;
        RECT 102.100 92.865 103.000 92.935 ;
        RECT 101.370 92.725 103.000 92.865 ;
        RECT 101.370 92.215 101.510 92.725 ;
        RECT 87.965 91.515 101.510 92.215 ;
        RECT 102.100 91.975 103.000 92.725 ;
        RECT 101.370 85.975 101.510 91.515 ;
        RECT 113.480 91.750 113.620 93.535 ;
        RECT 114.105 93.135 115.005 93.535 ;
        RECT 114.095 91.750 114.995 92.285 ;
        RECT 113.480 91.610 114.995 91.750 ;
        RECT 111.800 89.500 112.700 90.460 ;
        RECT 113.480 90.125 113.620 91.610 ;
        RECT 114.095 91.325 114.995 91.610 ;
        RECT 114.105 90.125 115.005 90.460 ;
        RECT 113.480 89.985 115.005 90.125 ;
        RECT 114.105 89.500 115.005 89.985 ;
        RECT 112.180 87.990 112.320 89.500 ;
        RECT 123.520 89.375 124.250 90.145 ;
        RECT 112.180 87.850 114.830 87.990 ;
        RECT 101.870 86.465 103.000 87.635 ;
        RECT 114.690 86.495 114.830 87.850 ;
        RECT 114.330 86.095 115.230 86.495 ;
        RECT 102.025 85.975 102.925 86.005 ;
        RECT 101.370 85.835 102.925 85.975 ;
        RECT 102.025 85.045 102.925 85.835 ;
        RECT 113.715 85.955 115.230 86.095 ;
        RECT 111.885 84.575 113.015 85.745 ;
        RECT 110.370 83.250 111.500 84.420 ;
        RECT 113.715 84.115 113.855 85.955 ;
        RECT 114.330 85.535 115.230 85.955 ;
        RECT 123.520 85.625 124.250 86.395 ;
        RECT 114.330 84.115 115.230 84.675 ;
        RECT 113.715 83.975 115.230 84.115 ;
        RECT 111.885 82.690 113.015 83.860 ;
        RECT 113.715 82.465 113.855 83.975 ;
        RECT 114.330 83.715 115.230 83.975 ;
        RECT 123.420 83.690 124.550 84.860 ;
        RECT 114.330 82.465 115.230 82.855 ;
        RECT 113.715 82.325 115.230 82.465 ;
        RECT 87.905 81.445 88.605 81.495 ;
        RECT 87.905 80.745 94.990 81.445 ;
        RECT 94.290 79.705 94.990 80.745 ;
        RECT 101.870 79.840 103.000 81.010 ;
        RECT 111.885 80.865 113.015 82.035 ;
        RECT 113.715 80.600 113.855 82.325 ;
        RECT 114.330 81.895 115.230 82.325 ;
        RECT 123.360 81.120 124.490 82.290 ;
        RECT 114.340 80.600 115.240 81.035 ;
        RECT 113.715 80.460 115.240 80.600 ;
        RECT 94.190 79.570 95.090 79.705 ;
        RECT 98.765 79.585 99.665 79.700 ;
        RECT 98.765 79.570 107.220 79.585 ;
        RECT 94.190 78.885 107.220 79.570 ;
        RECT 111.885 78.990 113.015 80.160 ;
        RECT 94.190 78.870 99.665 78.885 ;
        RECT 94.190 78.745 95.090 78.870 ;
        RECT 89.795 73.610 90.925 74.780 ;
        RECT 94.210 72.715 95.110 73.045 ;
        RECT 95.320 72.715 95.460 78.870 ;
        RECT 94.210 72.415 95.460 72.715 ;
        RECT 94.210 72.085 95.110 72.415 ;
        RECT 89.445 66.905 90.575 68.075 ;
        RECT 94.170 66.395 95.070 66.930 ;
        RECT 95.320 66.395 95.460 72.415 ;
        RECT 94.170 66.095 95.460 66.395 ;
        RECT 94.170 65.970 95.070 66.095 ;
        RECT 73.695 62.410 76.065 64.740 ;
        RECT 89.445 60.790 90.575 61.960 ;
        RECT 94.210 59.905 95.110 60.505 ;
        RECT 95.320 59.905 95.460 66.095 ;
        RECT 94.210 59.765 95.460 59.905 ;
        RECT 96.765 77.230 97.065 78.870 ;
        RECT 98.765 78.740 99.665 78.870 ;
        RECT 97.265 77.230 98.165 77.560 ;
        RECT 96.765 76.930 98.165 77.230 ;
        RECT 96.765 72.740 97.065 76.930 ;
        RECT 97.265 76.600 98.165 76.930 ;
        RECT 98.605 73.620 99.735 74.790 ;
        RECT 98.765 72.740 99.665 73.070 ;
        RECT 96.765 72.440 99.665 72.740 ;
        RECT 96.765 70.265 97.065 72.440 ;
        RECT 98.765 72.110 99.665 72.440 ;
        RECT 106.520 70.875 107.220 78.885 ;
        RECT 113.715 78.795 113.855 80.460 ;
        RECT 114.340 80.075 115.240 80.460 ;
        RECT 114.340 78.795 115.240 79.215 ;
        RECT 113.715 78.655 115.240 78.795 ;
        RECT 111.885 77.170 113.015 78.340 ;
        RECT 113.715 76.970 113.855 78.655 ;
        RECT 114.340 78.255 115.240 78.655 ;
        RECT 123.470 78.615 124.600 79.785 ;
        RECT 114.340 76.970 115.240 77.390 ;
        RECT 113.715 76.830 115.240 76.970 ;
        RECT 111.885 75.430 113.015 76.600 ;
        RECT 113.715 75.165 113.855 76.830 ;
        RECT 114.340 76.430 115.240 76.830 ;
        RECT 123.470 76.005 124.600 77.175 ;
        RECT 114.330 75.165 115.230 75.580 ;
        RECT 113.715 75.025 115.230 75.165 ;
        RECT 111.885 73.595 113.015 74.765 ;
        RECT 113.715 73.345 113.855 75.025 ;
        RECT 114.330 74.620 115.230 75.025 ;
        RECT 114.340 73.345 115.240 73.755 ;
        RECT 123.470 73.520 124.600 74.690 ;
        RECT 113.715 73.205 115.240 73.345 ;
        RECT 114.340 72.795 115.240 73.205 ;
        RECT 123.555 72.035 124.285 72.805 ;
        RECT 135.815 72.285 135.955 100.590 ;
        RECT 142.075 97.875 142.215 100.590 ;
        RECT 142.765 100.340 143.895 101.510 ;
        RECT 144.750 101.310 144.890 101.870 ;
        RECT 144.370 100.350 145.270 101.310 ;
        RECT 158.540 100.860 158.680 103.090 ;
        RECT 159.340 101.520 160.470 102.690 ;
        RECT 160.915 102.140 161.815 102.585 ;
        RECT 160.915 102.000 163.540 102.140 ;
        RECT 160.915 101.625 161.815 102.000 ;
        RECT 161.060 100.860 161.200 101.625 ;
        RECT 158.540 100.720 161.200 100.860 ;
        RECT 142.765 98.395 143.895 99.565 ;
        RECT 144.575 99.075 145.475 99.485 ;
        RECT 144.285 98.935 145.475 99.075 ;
        RECT 144.285 97.875 144.425 98.935 ;
        RECT 144.575 98.525 145.475 98.935 ;
        RECT 142.075 97.735 144.425 97.875 ;
        RECT 143.555 95.710 143.695 97.735 ;
        RECT 145.035 96.855 146.165 98.025 ;
        RECT 146.655 97.065 147.555 98.025 ;
        RECT 147.035 95.710 147.175 97.065 ;
        RECT 148.190 96.855 149.320 98.025 ;
        RECT 160.555 97.580 160.695 100.720 ;
        RECT 161.415 100.095 162.545 101.265 ;
        RECT 163.400 101.065 163.540 102.000 ;
        RECT 163.020 100.105 163.920 101.065 ;
        RECT 161.415 98.150 162.545 99.320 ;
        RECT 163.225 98.830 164.125 99.240 ;
        RECT 163.140 98.280 164.125 98.830 ;
        RECT 163.140 97.580 163.280 98.280 ;
        RECT 160.555 97.440 163.280 97.580 ;
        RECT 143.555 95.570 147.175 95.710 ;
        RECT 162.205 95.840 162.345 97.440 ;
        RECT 163.685 96.610 164.815 97.780 ;
        RECT 165.305 96.820 166.205 97.780 ;
        RECT 165.685 95.840 165.825 96.820 ;
        RECT 166.840 96.610 167.970 97.780 ;
        RECT 162.205 95.700 165.825 95.840 ;
        RECT 147.035 95.475 147.175 95.570 ;
        RECT 147.035 95.335 147.215 95.475 ;
        RECT 147.075 94.420 147.215 95.335 ;
        RECT 147.075 94.280 154.155 94.420 ;
        RECT 154.015 74.380 154.155 94.280 ;
        RECT 157.670 92.680 165.345 93.380 ;
        RECT 157.670 92.150 158.370 92.680 ;
        RECT 160.700 92.150 161.400 92.680 ;
        RECT 164.645 92.150 165.345 92.680 ;
        RECT 157.570 92.020 158.470 92.150 ;
        RECT 155.140 91.320 158.470 92.020 ;
        RECT 155.140 86.770 155.840 91.320 ;
        RECT 157.570 91.190 158.470 91.320 ;
        RECT 159.040 90.975 160.170 92.145 ;
        RECT 160.575 91.190 161.475 92.150 ;
        RECT 162.040 90.975 163.170 92.145 ;
        RECT 164.545 91.190 165.445 92.150 ;
        RECT 156.790 89.565 157.920 90.735 ;
        RECT 156.455 87.890 157.585 89.060 ;
        RECT 158.125 88.115 159.025 89.075 ;
        RECT 158.325 87.095 159.025 88.115 ;
        RECT 157.185 86.900 159.025 87.095 ;
        RECT 157.085 86.770 159.025 86.900 ;
        RECT 155.080 86.395 159.025 86.770 ;
        RECT 155.080 86.070 157.985 86.395 ;
        RECT 155.080 83.490 155.780 86.070 ;
        RECT 157.085 85.940 157.985 86.070 ;
        RECT 156.455 84.270 157.585 85.440 ;
        RECT 157.085 83.490 157.985 83.620 ;
        RECT 155.080 83.285 157.985 83.490 ;
        RECT 155.065 82.790 157.985 83.285 ;
        RECT 155.065 82.585 155.780 82.790 ;
        RECT 157.085 82.660 157.985 82.790 ;
        RECT 155.065 76.960 155.765 82.585 ;
        RECT 156.455 80.520 157.585 81.690 ;
        RECT 158.125 80.620 159.025 81.580 ;
        RECT 157.130 78.915 158.260 80.085 ;
        RECT 158.505 78.450 158.645 80.620 ;
        RECT 158.125 77.490 159.025 78.450 ;
        RECT 158.490 76.960 158.630 77.490 ;
        RECT 159.540 77.425 160.670 78.595 ;
        RECT 161.025 77.465 161.925 78.425 ;
        RECT 162.270 77.465 163.400 78.635 ;
        RECT 164.545 78.500 165.445 78.680 ;
        RECT 164.545 78.450 176.250 78.500 ;
        RECT 164.545 77.810 176.475 78.450 ;
        RECT 164.545 77.800 176.250 77.810 ;
        RECT 164.545 77.720 165.445 77.800 ;
        RECT 155.065 76.715 158.980 76.960 ;
        RECT 161.090 76.715 161.790 77.465 ;
        RECT 164.645 76.715 165.345 77.720 ;
        RECT 155.065 76.260 165.345 76.715 ;
        RECT 158.560 76.015 165.345 76.260 ;
        RECT 163.205 74.380 163.805 74.630 ;
        RECT 154.015 74.240 163.805 74.380 ;
        RECT 163.205 73.990 163.805 74.240 ;
        RECT 135.795 72.145 135.955 72.285 ;
        RECT 108.540 71.285 122.105 71.985 ;
        RECT 108.540 71.005 109.240 71.285 ;
        RECT 108.225 70.875 109.240 71.005 ;
        RECT 97.265 70.265 98.165 70.595 ;
        RECT 96.765 69.965 98.165 70.265 ;
        RECT 106.520 70.175 109.240 70.875 ;
        RECT 108.225 70.045 109.125 70.175 ;
        RECT 96.765 66.220 97.065 69.965 ;
        RECT 97.265 69.635 98.165 69.965 ;
        RECT 109.445 69.385 110.575 70.555 ;
        RECT 121.405 69.090 122.105 71.285 ;
        RECT 124.860 71.165 125.440 71.360 ;
        RECT 135.795 71.165 135.935 72.145 ;
        RECT 124.860 71.025 135.935 71.165 ;
        RECT 123.285 69.745 124.415 70.915 ;
        RECT 124.860 70.720 125.440 71.025 ;
        RECT 121.305 68.130 122.205 69.090 ;
        RECT 98.590 66.915 99.720 68.085 ;
        RECT 99.955 66.220 100.855 66.910 ;
        RECT 109.445 66.340 110.575 67.510 ;
        RECT 96.765 66.080 100.855 66.220 ;
        RECT 96.765 63.980 97.065 66.080 ;
        RECT 99.955 65.950 100.855 66.080 ;
        RECT 97.265 63.980 98.165 64.310 ;
        RECT 96.765 63.680 98.165 63.980 ;
        RECT 96.765 60.110 97.065 63.680 ;
        RECT 97.265 63.350 98.165 63.680 ;
        RECT 98.625 60.820 99.755 61.990 ;
        RECT 99.955 60.110 100.855 60.505 ;
        RECT 96.765 59.810 100.855 60.110 ;
        RECT 94.210 59.545 95.110 59.765 ;
        RECT 97.565 58.235 97.865 59.810 ;
        RECT 99.955 59.545 100.855 59.810 ;
        RECT 97.265 57.275 98.165 58.235 ;
        RECT 88.455 54.395 89.585 55.565 ;
        RECT 98.580 54.415 99.710 55.585 ;
        RECT 147.665 52.545 148.795 53.715 ;
        RECT 190.545 49.675 192.915 52.005 ;
        RECT 190.945 43.835 192.515 45.365 ;
        RECT 180.615 41.625 182.185 43.155 ;
        RECT 158.680 39.705 160.250 41.235 ;
        RECT 136.340 38.040 137.910 39.570 ;
        RECT 114.165 36.500 115.735 38.030 ;
      LAYER met3 ;
        RECT 150.115 248.675 150.415 248.680 ;
        RECT 149.900 247.905 150.630 248.675 ;
        RECT 158.095 248.045 158.825 248.815 ;
        RECT 150.115 244.505 150.415 247.905 ;
        RECT 158.310 244.505 158.610 248.045 ;
        RECT 150.115 244.205 158.610 244.505 ;
        RECT 150.115 241.500 150.415 244.205 ;
        RECT 158.310 241.735 158.610 244.205 ;
        RECT 149.900 240.730 150.630 241.500 ;
        RECT 158.095 240.965 158.825 241.735 ;
        RECT 150.115 234.550 150.415 240.730 ;
        RECT 158.310 234.865 158.610 240.965 ;
        RECT 149.900 233.780 150.630 234.550 ;
        RECT 158.095 234.095 158.825 234.865 ;
        RECT 150.115 227.525 150.415 233.780 ;
        RECT 158.310 227.525 158.610 234.095 ;
        RECT 148.130 227.240 148.860 227.475 ;
        RECT 149.900 227.240 150.630 227.525 ;
        RECT 148.130 226.940 150.630 227.240 ;
        RECT 148.130 226.705 148.860 226.940 ;
        RECT 149.900 226.755 150.630 226.940 ;
        RECT 158.095 226.755 158.825 227.525 ;
        RECT 105.545 225.095 106.675 225.595 ;
        RECT 105.545 224.795 109.820 225.095 ;
        RECT 105.545 224.425 106.675 224.795 ;
        RECT 109.520 223.295 109.820 224.795 ;
        RECT 149.900 223.725 150.630 224.495 ;
        RECT 150.115 223.295 150.415 223.725 ;
        RECT 109.520 222.995 150.415 223.295 ;
        RECT 158.310 208.460 158.610 226.755 ;
        RECT 158.065 207.690 158.795 208.460 ;
        RECT 158.310 201.670 158.610 207.690 ;
        RECT 158.065 200.900 158.795 201.670 ;
        RECT 69.985 183.655 72.365 183.815 ;
        RECT 73.695 183.655 76.065 183.820 ;
        RECT 69.985 181.655 76.065 183.655 ;
        RECT 69.985 181.495 72.365 181.655 ;
        RECT 73.695 181.490 76.065 181.655 ;
        RECT 190.545 182.670 192.915 182.835 ;
        RECT 196.075 182.670 198.455 182.830 ;
        RECT 190.545 180.670 198.455 182.670 ;
        RECT 190.545 180.505 192.915 180.670 ;
        RECT 196.075 180.510 198.455 180.670 ;
        RECT 123.965 143.730 124.695 143.850 ;
        RECT 94.605 143.715 124.695 143.730 ;
        RECT 93.255 143.430 124.695 143.715 ;
        RECT 93.255 143.415 94.905 143.430 ;
        RECT 93.255 136.510 93.555 143.415 ;
        RECT 123.965 143.080 124.695 143.430 ;
        RECT 96.275 136.510 97.405 137.260 ;
        RECT 93.255 136.210 97.405 136.510 ;
        RECT 93.255 126.640 93.555 136.210 ;
        RECT 96.275 136.090 97.405 136.210 ;
        RECT 105.260 136.125 106.390 137.295 ;
        RECT 105.675 134.620 105.975 136.125 ;
        RECT 115.755 136.065 116.885 137.235 ;
        RECT 115.940 135.045 116.240 136.065 ;
        RECT 104.010 134.320 105.975 134.620 ;
        RECT 114.375 134.745 116.320 135.045 ;
        RECT 96.275 126.640 97.405 127.350 ;
        RECT 93.255 126.340 97.405 126.640 ;
        RECT 96.275 126.180 97.405 126.340 ;
        RECT 104.010 127.060 104.310 134.320 ;
        RECT 105.260 127.060 106.390 127.385 ;
        RECT 104.010 126.760 106.390 127.060 ;
        RECT 96.275 116.545 97.405 117.195 ;
        RECT 95.310 116.245 97.405 116.545 ;
        RECT 95.310 107.635 95.610 116.245 ;
        RECT 96.275 116.025 97.405 116.245 ;
        RECT 104.010 116.935 104.310 126.760 ;
        RECT 105.260 126.215 106.390 126.760 ;
        RECT 114.375 126.780 114.675 134.745 ;
        RECT 172.500 132.895 173.230 132.930 ;
        RECT 155.250 132.195 173.230 132.895 ;
        RECT 146.945 130.365 148.075 130.560 ;
        RECT 145.255 129.665 148.075 130.365 ;
        RECT 145.255 128.835 145.955 129.665 ;
        RECT 146.945 129.390 148.075 129.665 ;
        RECT 145.040 128.610 146.170 128.835 ;
        RECT 143.920 127.910 146.170 128.610 ;
        RECT 155.250 128.150 155.950 132.195 ;
        RECT 172.500 132.160 173.230 132.195 ;
        RECT 165.275 130.365 166.405 130.560 ;
        RECT 163.585 129.665 166.405 130.365 ;
        RECT 163.585 128.835 164.285 129.665 ;
        RECT 165.275 129.390 166.405 129.665 ;
        RECT 163.370 128.610 164.500 128.835 ;
        RECT 115.755 126.780 116.885 127.340 ;
        RECT 143.920 127.270 144.620 127.910 ;
        RECT 145.040 127.665 146.170 127.910 ;
        RECT 143.920 127.255 145.140 127.270 ;
        RECT 114.375 126.480 116.885 126.780 ;
        RECT 105.260 116.935 106.390 117.370 ;
        RECT 104.010 116.635 106.390 116.935 ;
        RECT 102.830 110.790 103.560 111.025 ;
        RECT 104.010 110.790 104.310 116.635 ;
        RECT 105.260 116.200 106.390 116.635 ;
        RECT 114.375 117.030 114.675 126.480 ;
        RECT 115.755 126.170 116.885 126.480 ;
        RECT 141.875 126.555 145.140 127.255 ;
        RECT 155.075 126.980 156.205 128.150 ;
        RECT 162.335 127.910 164.500 128.610 ;
        RECT 162.335 127.340 163.035 127.910 ;
        RECT 163.370 127.665 164.500 127.910 ;
        RECT 160.205 127.270 163.255 127.340 ;
        RECT 141.875 125.765 142.575 126.555 ;
        RECT 144.010 126.100 145.140 126.555 ;
        RECT 160.205 126.640 163.470 127.270 ;
        RECT 160.205 125.765 160.905 126.640 ;
        RECT 162.340 126.100 163.470 126.640 ;
        RECT 141.660 125.385 142.790 125.765 ;
        RECT 159.990 125.470 161.120 125.765 ;
        RECT 138.705 124.685 142.790 125.385 ;
        RECT 138.705 123.605 139.405 124.685 ;
        RECT 141.660 124.595 142.790 124.685 ;
        RECT 157.035 124.770 161.120 125.470 ;
        RECT 157.035 123.625 157.735 124.770 ;
        RECT 159.990 124.595 161.120 124.770 ;
        RECT 138.445 122.435 139.575 123.605 ;
        RECT 156.775 122.455 157.905 123.625 ;
        RECT 138.720 120.850 139.420 122.435 ;
        RECT 140.980 120.850 142.110 121.225 ;
        RECT 138.720 120.150 142.110 120.850 ;
        RECT 157.050 120.990 157.750 122.455 ;
        RECT 159.310 120.990 160.440 121.225 ;
        RECT 157.050 120.290 160.440 120.990 ;
        RECT 140.980 120.055 142.110 120.150 ;
        RECT 159.310 120.055 160.440 120.290 ;
        RECT 141.335 119.075 142.035 120.055 ;
        RECT 143.055 119.075 144.185 119.800 ;
        RECT 141.335 118.630 144.185 119.075 ;
        RECT 159.665 119.215 160.365 120.055 ;
        RECT 161.385 119.215 162.515 119.800 ;
        RECT 159.665 118.630 162.515 119.215 ;
        RECT 141.335 118.375 143.970 118.630 ;
        RECT 159.665 118.515 162.300 118.630 ;
        RECT 143.270 117.855 143.970 118.375 ;
        RECT 161.600 117.855 162.300 118.515 ;
        RECT 115.755 117.030 116.885 117.485 ;
        RECT 124.800 117.235 125.930 117.635 ;
        RECT 114.375 116.730 116.885 117.030 ;
        RECT 102.830 110.490 104.310 110.790 ;
        RECT 102.830 110.255 103.560 110.490 ;
        RECT 96.275 107.755 97.405 108.190 ;
        RECT 104.010 108.055 104.310 110.490 ;
        RECT 105.260 108.065 106.390 108.165 ;
        RECT 114.375 108.065 114.675 116.730 ;
        RECT 115.755 116.315 116.885 116.730 ;
        RECT 123.250 116.935 125.930 117.235 ;
        RECT 115.755 108.065 116.885 108.310 ;
        RECT 105.260 108.055 116.885 108.065 ;
        RECT 104.010 107.765 116.885 108.055 ;
        RECT 104.010 107.755 106.390 107.765 ;
        RECT 96.275 107.635 104.310 107.755 ;
        RECT 95.310 107.455 104.310 107.635 ;
        RECT 95.310 107.335 97.405 107.455 ;
        RECT 96.275 107.020 97.405 107.335 ;
        RECT 105.260 106.995 106.390 107.755 ;
        RECT 115.755 107.140 116.885 107.765 ;
        RECT 123.250 107.545 123.550 116.935 ;
        RECT 124.800 116.465 125.930 116.935 ;
        RECT 143.055 116.685 144.185 117.855 ;
        RECT 161.385 116.685 162.515 117.855 ;
        RECT 143.135 115.940 143.835 116.685 ;
        RECT 145.325 115.940 146.455 116.315 ;
        RECT 143.135 115.240 146.455 115.940 ;
        RECT 145.325 115.145 146.455 115.240 ;
        RECT 148.480 115.960 149.610 116.315 ;
        RECT 161.465 115.960 162.165 116.685 ;
        RECT 163.655 115.960 164.785 116.315 ;
        RECT 148.480 115.260 164.785 115.960 ;
        RECT 148.480 115.145 149.610 115.260 ;
        RECT 145.540 114.820 146.240 115.145 ;
        RECT 148.705 114.820 149.405 115.145 ;
        RECT 145.540 114.120 149.405 114.820 ;
        RECT 146.705 112.075 147.835 112.270 ;
        RECT 144.965 111.375 147.835 112.075 ;
        RECT 144.965 110.545 145.665 111.375 ;
        RECT 146.705 111.100 147.835 111.375 ;
        RECT 144.750 110.320 145.880 110.545 ;
        RECT 143.735 109.620 145.880 110.320 ;
        RECT 143.735 109.110 144.435 109.620 ;
        RECT 144.750 109.375 145.880 109.620 ;
        RECT 141.390 108.980 144.440 109.110 ;
        RECT 141.390 108.410 144.850 108.980 ;
        RECT 124.395 107.545 125.525 108.010 ;
        RECT 123.250 107.245 125.525 107.545 ;
        RECT 141.390 107.475 142.090 108.410 ;
        RECT 143.720 107.810 144.850 108.410 ;
        RECT 123.250 106.695 123.550 107.245 ;
        RECT 124.395 106.840 125.525 107.245 ;
        RECT 141.370 107.240 142.500 107.475 ;
        RECT 100.980 106.395 123.550 106.695 ;
        RECT 138.220 106.540 142.500 107.240 ;
        RECT 100.980 100.555 101.280 106.395 ;
        RECT 108.935 104.130 109.235 106.395 ;
        RECT 138.220 105.335 138.920 106.540 ;
        RECT 141.370 106.305 142.500 106.540 ;
        RECT 138.155 104.165 139.285 105.335 ;
        RECT 108.750 103.360 109.480 104.130 ;
        RECT 138.220 102.470 138.920 104.165 ;
        RECT 140.690 102.470 141.820 102.935 ;
        RECT 138.220 101.770 141.820 102.470 ;
        RECT 140.690 101.765 141.820 101.770 ;
        RECT 101.870 100.555 103.000 100.990 ;
        RECT 100.980 100.255 103.000 100.555 ;
        RECT 98.310 93.815 99.040 94.095 ;
        RECT 100.980 93.815 101.280 100.255 ;
        RECT 101.870 99.820 103.000 100.255 ;
        RECT 141.045 100.695 141.745 101.765 ;
        RECT 142.765 100.695 143.895 101.510 ;
        RECT 141.045 100.340 143.895 100.695 ;
        RECT 141.045 99.995 143.680 100.340 ;
        RECT 142.980 99.565 143.680 99.995 ;
        RECT 142.765 98.395 143.895 99.565 ;
        RECT 142.845 97.560 143.545 98.395 ;
        RECT 145.035 97.560 146.165 98.025 ;
        RECT 142.845 96.860 146.165 97.560 ;
        RECT 145.035 96.855 146.165 96.860 ;
        RECT 148.190 97.325 149.320 98.025 ;
        RECT 153.810 97.325 154.510 115.260 ;
        RECT 163.655 115.145 164.785 115.260 ;
        RECT 166.810 115.145 167.940 116.315 ;
        RECT 164.000 114.840 164.700 115.145 ;
        RECT 167.025 114.840 167.725 115.145 ;
        RECT 164.000 114.140 167.725 114.840 ;
        RECT 165.305 111.830 166.435 112.025 ;
        RECT 163.615 111.130 166.435 111.830 ;
        RECT 163.615 110.300 164.315 111.130 ;
        RECT 165.305 110.855 166.435 111.130 ;
        RECT 163.400 110.075 164.530 110.300 ;
        RECT 162.360 109.375 164.530 110.075 ;
        RECT 162.360 108.865 163.060 109.375 ;
        RECT 163.400 109.130 164.530 109.375 ;
        RECT 160.020 108.735 163.070 108.865 ;
        RECT 160.020 108.165 163.500 108.735 ;
        RECT 160.020 107.230 160.720 108.165 ;
        RECT 162.360 108.150 163.500 108.165 ;
        RECT 162.370 107.565 163.500 108.150 ;
        RECT 160.020 106.995 161.150 107.230 ;
        RECT 156.850 106.295 161.150 106.995 ;
        RECT 156.850 105.105 157.550 106.295 ;
        RECT 160.020 106.060 161.150 106.295 ;
        RECT 156.805 103.935 157.935 105.105 ;
        RECT 156.850 102.455 157.550 103.935 ;
        RECT 159.340 102.455 160.470 102.690 ;
        RECT 156.850 101.755 160.470 102.455 ;
        RECT 159.340 101.520 160.470 101.755 ;
        RECT 159.695 100.680 160.395 101.520 ;
        RECT 161.415 100.680 162.545 101.265 ;
        RECT 159.695 100.095 162.545 100.680 ;
        RECT 159.695 99.980 162.330 100.095 ;
        RECT 161.630 99.320 162.330 99.980 ;
        RECT 161.415 98.150 162.545 99.320 ;
        RECT 161.495 97.325 162.195 98.150 ;
        RECT 163.685 97.325 164.815 97.780 ;
        RECT 148.190 96.855 164.815 97.325 ;
        RECT 145.250 96.440 145.950 96.855 ;
        RECT 148.405 96.625 164.815 96.855 ;
        RECT 148.405 96.440 149.115 96.625 ;
        RECT 145.250 95.740 149.115 96.440 ;
        RECT 152.920 95.960 153.620 96.625 ;
        RECT 163.685 96.610 164.815 96.625 ;
        RECT 166.840 96.610 167.970 97.780 ;
        RECT 163.900 96.205 164.600 96.610 ;
        RECT 167.065 96.205 167.765 96.610 ;
        RECT 152.920 95.220 153.695 95.960 ;
        RECT 163.900 95.505 167.765 96.205 ;
        RECT 152.975 95.180 153.695 95.220 ;
        RECT 101.870 93.815 103.000 94.300 ;
        RECT 98.310 93.515 103.000 93.815 ;
        RECT 98.310 93.325 99.040 93.515 ;
        RECT 101.870 93.130 103.000 93.515 ;
        RECT 155.685 93.930 160.355 93.960 ;
        RECT 155.685 93.260 162.955 93.930 ;
        RECT 155.685 90.515 156.385 93.260 ;
        RECT 159.275 93.230 162.955 93.260 ;
        RECT 159.275 92.145 159.975 93.230 ;
        RECT 162.255 92.145 162.955 93.230 ;
        RECT 159.040 90.975 160.170 92.145 ;
        RECT 162.040 90.975 163.170 92.145 ;
        RECT 156.790 90.515 157.920 90.735 ;
        RECT 123.325 89.170 124.445 90.350 ;
        RECT 154.490 89.815 157.920 90.515 ;
        RECT 154.490 88.625 155.190 89.815 ;
        RECT 156.790 89.565 157.920 89.815 ;
        RECT 156.455 88.625 157.585 89.060 ;
        RECT 154.490 88.325 157.585 88.625 ;
        RECT 101.870 87.200 103.000 87.635 ;
        RECT 100.970 86.900 103.000 87.200 ;
        RECT 100.970 80.720 101.270 86.900 ;
        RECT 101.870 86.465 103.000 86.900 ;
        RECT 111.885 84.575 113.015 85.745 ;
        RECT 123.325 85.420 124.445 86.600 ;
        RECT 154.490 85.585 155.190 88.325 ;
        RECT 156.455 87.890 157.585 88.325 ;
        RECT 154.490 85.005 155.255 85.585 ;
        RECT 156.455 85.005 157.585 85.440 ;
        RECT 154.490 84.885 157.585 85.005 ;
        RECT 110.370 83.250 111.500 84.420 ;
        RECT 112.300 83.860 112.600 84.575 ;
        RECT 110.910 81.705 111.210 83.250 ;
        RECT 111.885 82.690 113.015 83.860 ;
        RECT 123.420 83.690 124.550 84.860 ;
        RECT 154.550 84.705 157.585 84.885 ;
        RECT 112.300 82.035 112.600 82.690 ;
        RECT 123.885 82.290 124.185 83.690 ;
        RECT 111.885 81.705 113.015 82.035 ;
        RECT 110.910 81.405 113.015 81.705 ;
        RECT 101.870 80.810 103.000 81.010 ;
        RECT 110.910 80.810 111.210 81.405 ;
        RECT 111.885 80.865 113.015 81.405 ;
        RECT 123.360 81.120 124.490 82.290 ;
        RECT 101.870 80.720 111.210 80.810 ;
        RECT 100.970 80.510 111.210 80.720 ;
        RECT 100.970 80.420 103.000 80.510 ;
        RECT 101.870 79.840 103.000 80.420 ;
        RECT 112.300 80.160 112.600 80.865 ;
        RECT 111.885 78.990 113.015 80.160 ;
        RECT 123.885 79.785 124.185 81.120 ;
        RECT 154.550 79.850 155.250 84.705 ;
        RECT 156.455 84.270 157.585 84.705 ;
        RECT 156.455 81.455 157.585 81.690 ;
        RECT 156.110 80.520 157.585 81.455 ;
        RECT 156.110 79.850 156.810 80.520 ;
        RECT 157.130 79.850 158.260 80.085 ;
        RECT 112.300 78.340 112.600 78.990 ;
        RECT 123.470 78.615 124.600 79.785 ;
        RECT 154.550 79.150 158.260 79.850 ;
        RECT 111.885 77.170 113.015 78.340 ;
        RECT 123.885 77.175 124.185 78.615 ;
        RECT 112.300 76.600 112.600 77.170 ;
        RECT 111.885 75.430 113.015 76.600 ;
        RECT 123.470 76.005 124.600 77.175 ;
        RECT 156.110 76.765 156.810 79.150 ;
        RECT 157.130 78.915 158.260 79.150 ;
        RECT 159.540 77.425 160.670 78.595 ;
        RECT 162.270 77.465 163.400 78.635 ;
        RECT 156.110 76.465 156.950 76.765 ;
        RECT 87.405 74.345 89.045 74.375 ;
        RECT 89.795 74.345 90.925 74.780 ;
        RECT 98.605 74.355 99.735 74.790 ;
        RECT 112.300 74.765 112.600 75.430 ;
        RECT 87.405 74.045 90.925 74.345 ;
        RECT 87.405 67.875 87.705 74.045 ;
        RECT 89.795 73.610 90.925 74.045 ;
        RECT 96.430 74.055 99.735 74.355 ;
        RECT 89.445 67.875 90.575 68.075 ;
        RECT 87.405 67.575 90.575 67.875 ;
        RECT 69.985 64.575 72.365 64.735 ;
        RECT 73.695 64.575 76.065 64.740 ;
        RECT 69.985 62.575 76.065 64.575 ;
        RECT 69.985 62.415 72.365 62.575 ;
        RECT 73.695 62.410 76.065 62.575 ;
        RECT 87.405 61.655 87.705 67.575 ;
        RECT 89.445 66.905 90.575 67.575 ;
        RECT 96.430 67.660 96.730 74.055 ;
        RECT 98.605 73.620 99.735 74.055 ;
        RECT 111.885 73.595 113.015 74.765 ;
        RECT 123.885 74.690 124.185 76.005 ;
        RECT 156.450 75.875 156.750 76.465 ;
        RECT 159.755 75.875 160.455 77.425 ;
        RECT 162.470 75.875 163.170 77.465 ;
        RECT 147.775 75.175 163.170 75.875 ;
        RECT 123.470 73.520 124.600 74.690 ;
        RECT 123.885 72.805 124.185 73.520 ;
        RECT 123.555 72.035 124.285 72.805 ;
        RECT 109.445 70.120 110.575 70.555 ;
        RECT 123.285 70.120 124.415 70.915 ;
        RECT 106.630 69.820 124.415 70.120 ;
        RECT 98.590 67.715 99.720 68.085 ;
        RECT 106.630 67.715 106.930 69.820 ;
        RECT 109.445 69.385 110.575 69.820 ;
        RECT 123.285 69.745 124.415 69.820 ;
        RECT 96.430 67.650 97.615 67.660 ;
        RECT 98.590 67.650 106.930 67.715 ;
        RECT 96.430 67.415 106.930 67.650 ;
        RECT 96.430 67.350 99.720 67.415 ;
        RECT 89.445 61.655 90.575 61.960 ;
        RECT 87.405 61.355 90.575 61.655 ;
        RECT 87.405 55.130 87.705 61.355 ;
        RECT 89.445 60.790 90.575 61.355 ;
        RECT 96.430 61.625 96.730 67.350 ;
        RECT 98.590 66.915 99.720 67.350 ;
        RECT 108.260 67.075 108.980 67.200 ;
        RECT 109.445 67.075 110.575 67.510 ;
        RECT 108.260 66.775 110.575 67.075 ;
        RECT 108.260 66.420 108.980 66.775 ;
        RECT 109.445 66.340 110.575 66.775 ;
        RECT 98.625 61.625 99.755 61.990 ;
        RECT 96.430 61.325 99.755 61.625 ;
        RECT 88.455 55.130 89.585 55.565 ;
        RECT 87.405 55.045 89.585 55.130 ;
        RECT 96.430 55.045 96.730 61.325 ;
        RECT 97.360 61.305 97.660 61.325 ;
        RECT 98.625 60.820 99.755 61.325 ;
        RECT 98.580 55.045 99.710 55.585 ;
        RECT 87.405 54.830 99.710 55.045 ;
        RECT 88.455 54.745 99.710 54.830 ;
        RECT 88.455 54.395 89.585 54.745 ;
        RECT 98.580 54.415 99.710 54.745 ;
        RECT 147.775 53.715 148.475 75.175 ;
        RECT 147.665 53.480 148.795 53.715 ;
        RECT 152.465 53.480 174.920 69.780 ;
        RECT 147.665 52.780 174.920 53.480 ;
        RECT 147.665 52.545 148.795 52.780 ;
        RECT 152.465 47.330 174.920 52.780 ;
        RECT 190.545 51.840 192.915 52.005 ;
        RECT 196.075 51.840 198.455 52.000 ;
        RECT 190.545 49.840 198.455 51.840 ;
        RECT 190.545 49.675 192.915 49.840 ;
        RECT 196.075 49.680 198.455 49.840 ;
        RECT 191.730 45.365 197.305 45.600 ;
        RECT 190.945 45.360 197.305 45.365 ;
        RECT 190.945 43.840 198.055 45.360 ;
        RECT 190.945 43.835 197.305 43.840 ;
        RECT 191.730 43.600 197.305 43.835 ;
        RECT 180.615 43.150 186.975 43.390 ;
        RECT 180.615 41.630 187.725 43.150 ;
        RECT 158.680 41.230 165.040 41.470 ;
        RECT 180.615 41.390 186.975 41.630 ;
        RECT 136.340 39.565 142.700 39.805 ;
        RECT 158.680 39.710 165.790 41.230 ;
        RECT 119.695 38.040 121.275 38.060 ;
        RECT 114.165 37.040 121.275 38.040 ;
        RECT 136.340 38.045 143.450 39.565 ;
        RECT 158.680 39.470 165.040 39.710 ;
        RECT 136.340 37.805 142.700 38.045 ;
        RECT 114.165 36.500 115.735 37.040 ;
        RECT 119.695 36.540 121.275 37.040 ;
      LAYER met4 ;
        RECT 56.355 260.075 56.655 260.780 ;
        RECT 60.035 260.075 60.335 260.780 ;
        RECT 63.715 260.075 64.015 260.780 ;
        RECT 67.395 260.075 67.695 260.780 ;
        RECT 71.075 260.075 71.375 260.780 ;
        RECT 74.755 260.075 75.055 260.780 ;
        RECT 78.435 260.075 78.735 260.780 ;
        RECT 82.115 260.075 82.415 260.780 ;
        RECT 85.795 260.075 86.095 260.780 ;
        RECT 89.475 260.075 89.775 260.780 ;
        RECT 93.155 260.075 93.455 260.780 ;
        RECT 96.835 260.075 97.135 260.780 ;
        RECT 100.515 260.075 100.815 260.780 ;
        RECT 104.195 260.075 104.495 260.780 ;
        RECT 107.875 260.075 108.175 260.780 ;
        RECT 111.555 260.075 111.855 260.780 ;
        RECT 115.235 260.075 115.535 260.780 ;
        RECT 118.915 260.075 119.215 260.780 ;
        RECT 122.595 260.075 122.895 260.780 ;
        RECT 126.275 260.075 126.575 260.780 ;
        RECT 129.955 260.075 130.255 260.780 ;
        RECT 133.635 260.075 133.935 260.780 ;
        RECT 137.315 260.075 137.615 260.780 ;
        RECT 140.995 260.075 141.295 260.780 ;
        RECT 55.855 259.780 141.295 260.075 ;
        RECT 144.675 259.780 144.975 260.780 ;
        RECT 148.355 259.780 148.655 260.780 ;
        RECT 152.035 259.780 152.335 260.780 ;
        RECT 155.715 259.780 156.015 260.780 ;
        RECT 159.395 259.780 159.695 260.780 ;
        RECT 163.075 259.780 163.375 260.780 ;
        RECT 166.755 259.780 167.055 260.780 ;
        RECT 170.435 259.780 170.735 260.780 ;
        RECT 174.115 259.780 174.415 260.780 ;
        RECT 177.795 259.780 178.095 260.780 ;
        RECT 181.475 259.780 181.775 260.780 ;
        RECT 185.155 259.780 185.455 260.780 ;
        RECT 188.835 259.780 189.135 260.780 ;
        RECT 192.515 259.780 192.815 260.780 ;
        RECT 196.195 259.780 196.495 260.780 ;
        RECT 199.875 259.780 200.175 260.780 ;
        RECT 203.555 259.780 203.855 260.780 ;
        RECT 207.235 259.780 207.535 260.780 ;
        RECT 210.915 259.780 211.215 260.780 ;
        RECT 55.855 259.775 141.135 259.780 ;
        RECT 55.855 183.675 57.855 259.775 ;
        RECT 70.010 183.675 72.340 183.820 ;
        RECT 55.855 181.675 72.450 183.675 ;
        RECT 196.100 182.690 198.430 182.835 ;
        RECT 210.720 182.690 212.720 259.170 ;
        RECT 55.855 64.595 57.855 181.675 ;
        RECT 70.010 181.490 72.340 181.675 ;
        RECT 196.100 180.690 212.720 182.690 ;
        RECT 196.100 180.505 198.430 180.690 ;
        RECT 152.970 95.205 153.700 95.935 ;
        RECT 123.320 89.195 124.450 90.325 ;
        RECT 123.735 87.290 124.035 89.195 ;
        RECT 109.935 86.990 124.035 87.290 ;
        RECT 109.935 78.765 110.235 86.990 ;
        RECT 123.735 86.575 124.035 86.990 ;
        RECT 123.320 85.445 124.450 86.575 ;
        RECT 108.315 78.745 110.235 78.765 ;
        RECT 107.300 78.465 110.235 78.745 ;
        RECT 107.300 78.445 108.615 78.465 ;
        RECT 107.300 66.960 107.600 78.445 ;
        RECT 152.985 69.640 153.685 95.205 ;
        RECT 108.255 66.960 108.985 67.175 ;
        RECT 107.300 66.660 108.985 66.960 ;
        RECT 108.255 66.445 108.985 66.660 ;
        RECT 70.010 64.595 72.340 64.740 ;
        RECT 55.855 62.595 72.450 64.595 ;
        RECT 55.855 54.285 57.855 62.595 ;
        RECT 70.010 62.410 72.340 62.595 ;
        RECT 55.855 54.275 57.065 54.285 ;
        RECT 57.075 54.275 57.855 54.285 ;
        RECT 55.855 36.025 57.855 54.275 ;
        RECT 152.605 47.470 174.780 69.640 ;
        RECT 196.100 51.860 198.430 52.005 ;
        RECT 210.720 51.860 212.720 180.690 ;
        RECT 196.100 49.860 212.720 51.860 ;
        RECT 196.100 49.675 198.430 49.860 ;
        RECT 197.265 45.365 210.100 45.600 ;
        RECT 196.500 43.835 210.100 45.365 ;
        RECT 197.265 43.600 210.100 43.835 ;
        RECT 186.170 41.625 187.700 43.155 ;
        RECT 164.235 39.705 165.765 41.235 ;
        RECT 141.895 39.300 143.425 39.570 ;
        RECT 119.720 37.970 121.250 38.065 ;
        RECT 141.895 38.040 143.525 39.300 ;
        RECT 119.720 36.535 121.380 37.970 ;
        RECT 54.365 35.020 54.965 36.020 ;
        RECT 76.445 35.020 77.045 36.020 ;
        RECT 98.525 35.020 99.125 36.020 ;
        RECT 120.380 35.690 121.380 36.535 ;
        RECT 142.525 35.850 143.525 38.040 ;
        RECT 120.605 35.020 121.205 35.690 ;
        RECT 142.685 35.020 143.285 35.850 ;
        RECT 164.505 35.515 165.505 39.705 ;
        RECT 186.655 35.810 187.655 41.625 ;
        RECT 164.765 35.020 165.365 35.515 ;
        RECT 186.845 35.020 187.445 35.810 ;
        RECT 208.100 35.690 210.100 43.600 ;
        RECT 210.720 43.995 212.720 49.860 ;
        RECT 210.720 43.985 211.645 43.995 ;
        RECT 211.655 43.985 212.720 43.995 ;
        RECT 210.720 36.025 212.720 43.985 ;
        RECT 208.925 35.020 209.525 35.690 ;
  END
END tt_um_Burrows_Katie
END LIBRARY

